-- code generated from the following source code:
--   ../rvm.ecl
--
-- with the following command:
--
--    ./eclat -notyB ../rvm.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 31);
       signal result : out value(0 to 1));
       
end entity;
architecture rtl of main is

  type t_state is (compute3364, \$10694_forever290\);
  signal state: t_state;
  type t_state_var7021 is (compute3367, \$10704_forever290\, \$10778_run286\, \$10801_forever3163135\, \$10805_forever3163133\, \$10859_forever3163136\, \$10863_forever3163133\, \$10872_forever3163137\, \$10876_forever3163133\, \$10885_forever3163138\, \$10889_forever3163133\, \$10905_forever3163139\, \$10909_forever3163133\, \$10932_forever3163140\, \$10936_forever3163133\, \$10945_forever3163141\, \$10949_forever3163133\, \$10958_forever3163142\, \$10962_forever3163133\, \$10971_forever3163143\, \$10975_forever3163133\, \$10998_forever3163144\, \$11002_forever3163133\, \$11011_forever3163145\, \$11015_forever3163133\, \$11024_forever3163146\, \$11028_forever3163133\, \$11036_loop3073149\, \$11057_forever3163147\, \$11061_forever3163133\, \$11073_forever3163148\, \$11077_forever3163133\, \$11090_forever3163150\, \$11094_forever3163133\, \$11113_forever3163151\, \$11117_forever3163133\, \$11126_forever3163152\, \$11130_forever3163133\, \$11139_forever3163153\, \$11143_forever3163133\, \$11164_forever3163154\, \$11168_forever3163133\, \$11177_forever3163155\, \$11181_forever3163133\, \$11196_loop2913158\, \$11244_forever3163156\, \$11248_forever3163133\, \$11259_forever3163157\, \$11263_forever3163133\, \$11272_forever3163159\, \$11276_forever3163133\, \$11285_forever3163160\, \$11289_forever3163133\, \$11311_forever3163161\, \$11315_forever3163133\, \$11343_forever3163162\, \$11347_forever3163133\, \$11356_forever3163163\, \$11360_forever3163133\, \$11370_forever3163164\, \$11374_forever3163133\, \$11398_forever3163165\, \$11402_forever3163133\, \$11412_forever3163166\, \$11416_forever3163133\, \$11425_forever3163167\, \$11429_forever3163133\, \$11437_loop3073170\, \$11458_forever3163168\, \$11462_forever3163133\, \$11474_forever3163169\, \$11478_forever3163133\, \$11496_forever3163171\, \$11500_forever3163133\, \$11510_forever3163172\, \$11514_forever3163133\, \$11525_forever3163173\, \$11529_forever3163133\, \$11584_forever3163174\, \$11588_forever3163133\, \$11604_forever3163175\, \$11608_forever3163133\, \$11619_forever3163176\, \$11623_forever3163133\, \$11633_forever3163177\, \$11637_forever3163133\, \$11647_forever3163178\, \$11651_forever3163133\, \$11683_forever3163179\, \$11687_forever3163133\, \$11698_forever3163180\, \$11702_forever3163133\, \$11720_forever3163181\, \$11724_forever3163133\, \$11764_forever3163182\, \$11768_forever3163133\, \$11779_forever3163183\, \$11783_forever3163133\, \$11793_forever3163184\, \$11797_forever3163133\, \$11834_forever3163185\, \$11838_forever3163133\, \$11867_forever3163186\, \$11871_forever3163133\, \$11881_forever3163187\, \$11885_forever3163133\, \$11895_forever3163188\, \$11899_forever3163133\, \$11933_forever3163189\, \$11937_forever3163133\, \$11951_forever3163190\, \$11955_forever3163133\, \$11992_forever3163191\, \$11996_forever3163133\, \$12006_forever3163192\, \$12010_forever3163133\, \$12020_forever3163193\, \$12024_forever3163133\, \$12061_forever3163194\, \$12065_forever3163133\, \$12075_forever3163195\, \$12079_forever3163133\, \$12089_forever3163196\, \$12093_forever3163133\, \$12130_forever3163197\, \$12134_forever3163133\, \$12144_forever3163198\, \$12148_forever3163133\, \$12158_forever3163199\, \$12162_forever3163133\, \$12203_forever3163200\, \$12207_forever3163133\, \$12217_forever3163201\, \$12221_forever3163133\, \$12240_forever3163202\, \$12244_forever3163133\, \$12253_forever3163203\, \$12257_forever3163133\, \$12267_forever3163204\, \$12271_forever3163133\, \$12281_forever3163205\, \$12285_forever3163133\, \$12326_forever3163206\, \$12330_forever3163133\, \$12340_forever3163207\, \$12344_forever3163133\, \$12363_forever3163208\, \$12367_forever3163133\, \$12376_forever3163209\, \$12380_forever3163133\, \$12390_forever3163210\, \$12394_forever3163133\, \$12404_forever3163211\, \$12408_forever3163133\, \$12449_forever3163212\, \$12453_forever3163133\, \$12463_forever3163213\, \$12467_forever3163133\, \$12486_forever3163214\, \$12490_forever3163133\, \$12499_forever3163215\, \$12503_forever3163133\, \$12513_forever3163216\, \$12517_forever3163133\, \$12527_forever3163217\, \$12531_forever3163133\, \$12573_forever3163218\, \$12577_forever3163133\, \$12621_forever3163219\, \$12625_forever3163133\, \$12634_forever3163220\, \$12638_forever3163133\, \$12648_forever3163221\, \$12652_forever3163133\, \$12662_forever3163222\, \$12666_forever3163133\, \$12707_forever3163223\, \$12711_forever3163133\, \$12723_forever3163225\, \$12727_forever3163133\, \$12734_forever3163224\, \$12738_forever3163133\, \$12747_forever3163226\, \$12751_forever3163133\, \$12761_forever3163227\, \$12765_forever3163133\, \$12806_forever3163228\, \$12810_forever3163133\, \$12820_forever3163229\, \$12824_forever3163133\, \$12834_forever3163230\, \$12838_forever3163133\, \$12847_forever3163231\, \$12851_forever3163133\, \$12861_forever3163232\, \$12865_forever3163133\, \$12906_forever3163233\, \$12910_forever3163133\, \$12920_forever3163234\, \$12924_forever3163133\, \$12934_forever3163235\, \$12938_forever3163133\, \$12947_forever3163236\, \$12951_forever3163133\, \$12961_forever3163237\, \$12965_forever3163133\, \$13006_forever3163238\, \$13010_forever3163133\, \$13020_forever3163239\, \$13024_forever3163133\, \$13034_forever3163240\, \$13038_forever3163133\, \$13047_forever3163241\, \$13051_forever3163133\, \$13061_forever3163242\, \$13065_forever3163133\, \$13106_forever3163243\, \$13110_forever3163133\, \$13120_forever3163244\, \$13124_forever3163133\, \$13134_forever3163245\, \$13138_forever3163133\, \$13147_forever3163246\, \$13151_forever3163133\, \$13161_forever3163247\, \$13165_forever3163133\, \$13194_forever3163248\, \$13198_forever3163133\, \$13206_forever3163249\, \$13210_forever3163133\, \$13242_forever3163250\, \$13246_forever3163133\, \$13257_forever3163251\, \$13261_forever3163133\, \$13270_forever3163252\, \$13274_forever3163133\, \$13283_forever3163253\, \$13287_forever3163133\, \$13305_forever3163254\, \$13309_forever3163133\, \$13318_list_tail2653256\, \$13339_forever3163255\, \$13343_forever3163133\, \$13360_forever3163257\, \$13364_forever3163133\, \$13374_forever3163258\, \$13378_forever3163133\, \$13388_forever3163259\, \$13392_forever3163133\, \$13420_forever3163260\, \$13424_forever3163133\, \$13434_forever3163261\, \$13438_forever3163133\, \$13451_forever3163262\, \$13455_forever3163133\, \$13474_forever3163263\, \$13478_forever3163133\, \$13487_forever3163264\, \$13491_forever3163133\, \$13500_list_tail2653266\, \$13521_forever3163265\, \$13525_forever3163133\, \$13537_forever3163267\, \$13541_forever3163133\, \$13560_forever3163268\, \$13564_forever3163133\, \$13573_forever3163269\, \$13577_forever3163133\, \$13587_forever3163270\, \$13591_forever3163133\, \$13618_forever3163271\, \$13622_forever3163133\, \$13632_forever3163272\, \$13636_forever3163133\, \$13653_forever3163273\, \$13657_forever3163133\, \$13676_forever3163274\, \$13680_forever3163133\, \$13689_list_tail2653276\, \$13710_forever3163275\, \$13714_forever3163133\, \$13731_forever3163277\, \$13735_forever3163133\, \$13761_forever3163278\, \$13765_forever3163133\, \$13775_forever3163279\, \$13779_forever3163133\, \$13796_forever3163280\, \$13800_forever3163133\, \$13821_forever3163281\, \$13825_forever3163133\, \$13842_forever3163282\, \$13846_forever3163133\, \$13856_forever3163283\, \$13860_forever3163133\, \$13878_forever3163284\, \$13882_forever3163133\, \$13892_forever3163134\, \$13896_forever3163133\, \$13905_forever3163285\, \$13909_forever3163133\, \$13931_forever3163286\, \$13935_forever3163133\, \$13950_forever3163287\, \$13954_forever3163133\, \$13977_forever3163288\, \$13981_forever3163133\, \$13991_forever3163289\, \$13995_forever3163133\, \$14004_forever3163290\, \$14008_forever3163133\, \$14037_forever3163291\, \$14041_forever3163133\, \$14050_forever3163292\, \$14054_forever3163133\, \$14064_forever3163293\, \$14068_forever3163133\, \$14090_forever3163294\, \$14094_forever3163133\, \$14104_forever3163295\, \$14108_forever3163133\, \$14117_forever3163296\, \$14121_forever3163133\, \$14150_forever3163297\, \$14154_forever3163133\, \$14163_forever3163298\, \$14167_forever3163133\, \$14177_forever3163299\, \$14181_forever3163133\, \$14203_forever3163300\, \$14207_forever3163133\, \$14217_forever3163301\, \$14221_forever3163133\, \$14230_forever3163302\, \$14234_forever3163133\, \$14263_forever3163303\, \$14267_forever3163133\, \$14276_forever3163304\, \$14280_forever3163133\, \$14290_forever3163305\, \$14294_forever3163133\, \$14311_forever3163306\, \$14315_forever3163133\, \$14325_forever3163307\, \$14329_forever3163133\, \$14338_forever3163308\, \$14342_forever3163133\, \$14369_forever3163309\, \$14373_forever3163133\, \$14382_forever3163310\, \$14386_forever3163133\, \$14396_forever3163311\, \$14400_forever3163133\, \$14423_forever3163312\, \$14427_forever3163133\, \$14437_forever3163313\, \$14441_forever3163133\, \$14450_forever3163314\, \$14454_forever3163133\, \$14464_forever3163315\, \$14468_forever3163133\, \$14481_decode_loop310\, \$14511_loop311\, \$14548_forever3163316\, \$14552_forever3163133\, \$14572_forever3163317\, \$14576_forever3163133\, \$14586_forever3163318\, \$14590_forever3163133\, \$14617_forever3163319\, \$14621_forever3163133\, \$14632_forever3163320\, \$14636_forever3163133\, \$14673_forever3163321\, \$14677_forever3163133\, \$14697_forever3163322\, \$14701_forever3163133\, \$14711_forever3163323\, \$14715_forever3163133\, \$14740_forever3163324\, \$14744_forever3163133\, \$14755_forever3163325\, \$14759_forever3163133\, \$14785_forever3163326\, \$14789_forever3163133\, \$14811_forever3163327\, \$14815_forever3163133\, \$14826_forever3163328\, \$14830_forever3163133\, \$14850_forever3163329\, \$14854_forever3163133\, \$14863_list_tail2653331\, \$14884_forever3163330\, \$14888_forever3163133\, \$14897_get_int268\, \$14939_get_int268\, \$14983_forever3163332\, \$14987_forever3163133\, \$14996_list_tail2653334\, \$15017_forever3163333\, \$15021_forever3163133\, \$15051_forever3163335\, \$15055_forever3163133\, \$15082_forever3163336\, \$15086_forever3163133\, \$15106_forever3163337\, \$15110_forever3163133\, \$15120_forever3163338\, \$15124_forever3163133\, \$15149_forever3163339\, \$15153_forever3163133\, \$15164_forever3163340\, \$15168_forever3163133\, \$15178_forever3163341\, \$15182_forever3163133\, \$15217_loop1312\, \$15240_loop23133355\, \$15282_forever3163342\, \$15286_forever3163133\, \$15332_forever3163343\, \$15336_forever3163133\, \$15355_forever3163344\, \$15359_forever3163133\, \$15378_forever3163345\, \$15382_forever3163133\, \$15391_len_aux3143348\, \$15413_forever3163346\, \$15417_forever3163133\, \$15439_forever3163347\, \$15443_forever3163133\, \$15496_forever3163349\, \$15500_forever3163133\, \$15519_forever3163350\, \$15523_forever3163133\, \$15542_forever3163351\, \$15546_forever3163133\, \$15555_len_aux3143354\, \$15577_forever3163352\, \$15581_forever3163133\, \$15603_forever3163353\, \$15607_forever3163133\, \$15663_forever3163356\, \$15667_forever3163133\, \$15686_forever3163357\, \$15690_forever3163133\, \$15710_forever3163358\, \$15714_forever3163133\, \$15724_len_aux3143361\, \$15746_forever3163359\, \$15750_forever3163133\, \$15772_forever3163360\, \$15776_forever3163133\, \$15788_get_int268\, pause_getI3378, pause_getI3397, pause_getI3404, pause_getI3418, pause_getI3425, pause_getI3433, pause_getI3443, pause_getI3450, pause_getI3459, pause_getI3471, pause_getI3478, pause_getI3487, pause_getI3494, pause_getI3505, pause_getI3511, pause_getI3519, pause_getI3528, pause_getI3536, pause_getI3540, pause_getI3548, pause_getI3553, pause_getI3557, pause_getI3568, pause_getI3572, pause_getI3581, pause_getI3587, pause_getI3597, pause_getI3605, pause_getI3609, pause_getI3617, pause_getI3622, pause_getI3626, pause_getI3638, pause_getI3644, pause_getI3656, pause_getI3668, pause_getI3675, pause_getI3684, pause_getI3690, pause_getI3695, pause_getI3706, pause_getI3712, pause_getI3725, pause_getI3733, pause_getI3737, pause_getI3741, pause_getI3749, pause_getI3754, pause_getI3758, pause_getI3762, pause_getI3770, pause_getI3778, pause_getI3782, pause_getI3790, pause_getI3795, pause_getI3799, pause_getI3810, pause_getI3814, pause_getI3825, pause_getI3829, pause_getI3840, pause_getI3844, pause_getI3853, pause_getI3861, pause_getI3865, pause_getI3869, pause_getI3877, pause_getI3882, pause_getI3886, pause_getI3897, pause_getI3901, pause_getI3912, pause_getI3916, pause_getI3925, pause_getI3933, pause_getI3937, pause_getI3941, pause_getI3949, pause_getI3954, pause_getI3958, pause_getI3969, pause_getI3973, pause_getI3984, pause_getI3988, pause_getI3997, pause_getI4005, pause_getI4009, pause_getI4013, pause_getI4021, pause_getI4026, pause_getI4030, pause_getI4034, pause_getI4043, pause_getI4051, pause_getI4055, pause_getI4063, pause_getI4068, pause_getI4072, pause_getI4076, pause_getI4081, pause_getI4094, pause_getI4098, pause_getI4109, pause_getI4117, pause_getI4121, pause_getI4125, pause_getI4133, pause_getI4138, pause_getI4142, pause_getI4156, pause_getI4160, pause_getI4169, pause_getI4177, pause_getI4181, pause_getI4185, pause_getI4193, pause_getI4198, pause_getI4202, pause_getI4207, pause_getI4220, pause_getI4224, pause_getI4233, pause_getI4241, pause_getI4245, pause_getI4249, pause_getI4257, pause_getI4262, pause_getI4266, pause_getI4271, pause_getI4284, pause_getI4288, pause_getI4297, pause_getI4305, pause_getI4309, pause_getI4313, pause_getI4321, pause_getI4326, pause_getI4330, pause_getI4335, pause_getI4348, pause_getI4352, pause_getI4361, pause_getI4369, pause_getI4373, pause_getI4377, pause_getI4385, pause_getI4390, pause_getI4394, pause_getI4404, pause_getI4411, pause_getI4426, pause_getI4430, pause_getI4441, pause_getI4445, pause_getI4454, pause_getI4462, pause_getI4466, pause_getI4470, pause_getI4478, pause_getI4483, pause_getI4487, pause_getI4497, pause_getI4504, pause_getI4519, pause_getI4523, pause_getI4534, pause_getI4538, pause_getI4547, pause_getI4555, pause_getI4559, pause_getI4563, pause_getI4571, pause_getI4576, pause_getI4580, pause_getI4590, pause_getI4597, pause_getI4612, pause_getI4616, pause_getI4627, pause_getI4631, pause_getI4642, pause_getI4650, pause_getI4654, pause_getI4658, pause_getI4666, pause_getI4671, pause_getI4675, pause_getI4714, pause_getI4721, pause_getI4738, pause_getI4742, pause_getI4753, pause_getI4757, pause_getI4766, pause_getI4774, pause_getI4778, pause_getI4782, pause_getI4790, pause_getI4795, pause_getI4799, pause_getI4818, pause_getI4822, pause_getI4833, pause_getI4837, pause_getI4846, pause_getI4854, pause_getI4858, pause_getI4862, pause_getI4870, pause_getI4875, pause_getI4879, pause_getI4897, pause_getI4901, pause_getI4912, pause_getI4916, pause_getI4925, pause_getI4933, pause_getI4937, pause_getI4941, pause_getI4949, pause_getI4954, pause_getI4958, pause_getI4976, pause_getI4980, pause_getI4991, pause_getI4995, pause_getI5004, pause_getI5012, pause_getI5016, pause_getI5020, pause_getI5028, pause_getI5033, pause_getI5037, pause_getI5055, pause_getI5059, pause_getI5070, pause_getI5074, pause_getI5083, pause_getI5091, pause_getI5095, pause_getI5099, pause_getI5107, pause_getI5112, pause_getI5116, pause_getI5134, pause_getI5138, pause_getI5149, pause_getI5153, pause_getI5162, pause_getI5170, pause_getI5174, pause_getI5178, pause_getI5186, pause_getI5191, pause_getI5195, pause_getI5204, pause_getI5212, pause_getI5216, pause_getI5220, pause_getI5228, pause_getI5233, pause_getI5237, pause_getI5251, pause_getI5255, pause_getI5263, pause_getI5271, pause_getI5278, pause_getI5285, pause_getI5290, pause_getI5299, pause_getI5305, pause_getI5310, pause_getI5314, pause_getI5326, pause_getI5332, pause_getI5343, pause_getI5350, pause_getI5359, pause_getI5366, pause_getI5376, pause_getI5383, pause_getI5400, pause_getI5404, pause_getI5416, pause_getI5422, pause_getI5431, pause_getI5439, pause_getI5443, pause_getI5447, pause_getI5455, pause_getI5460, pause_getI5464, pause_getI5470, pause_getI5477, pause_getI5484, pause_getI5489, pause_getI5505, pause_getI5511, pause_getI5520, pause_getI5528, pause_getI5532, pause_getI5536, pause_getI5544, pause_getI5549, pause_getI5553, pause_getI5565, pause_getI5571, pause_getI5601, pause_getI5605, pause_getI5613, pause_getI5619, pause_getI5640, pause_getI5644, pause_getI5652, pause_getI5657, pause_getI5661, pause_getI5665, pause_getI5669, pause_getI5677, pause_getI5682, pause_getI5686, pause_getI5698, pause_getI5704, pause_getI5715, pause_getI5722, pause_getI5731, pause_getI5737, pause_getI5749, pause_getI5755, pause_getI5766, pause_getI5773, pause_getI5782, pause_getI5788, pause_getI5800, pause_getI5806, pause_getI5817, pause_getI5824, pause_getI5833, pause_getI5839, pause_getI5851, pause_getI5857, pause_getI5867, pause_getI5874, pause_getI5883, pause_getI5889, pause_getI5893, pause_getI5903, pause_getI5911, pause_getI5915, pause_getI5923, pause_getI5928, pause_getI5932, pause_getI5936, pause_getI5948, pause_getI5955, pause_getI5961, pause_getI5971, pause_getI5978, pause_getI5986, pause_getI5995, pause_getI6003, pause_getI6007, pause_getI6015, pause_getI6020, pause_getI6024, pause_getI6029, pause_getI6035, pause_getI6046, pause_getI6050, pause_getI6060, pause_getI6067, pause_getI6075, pause_getI6084, pause_getI6092, pause_getI6096, pause_getI6104, pause_getI6109, pause_getI6113, pause_getI6118, pause_getI6124, pause_getI6132, pause_getI6136, pause_getI6146, pause_getI6154, pause_getI6158, pause_getI6166, pause_getI6171, pause_getI6175, pause_getI6179, pause_getI6188, pause_getI6196, pause_getI6200, pause_getI6208, pause_getI6213, pause_getI6217, pause_getI6228, pause_getI6232, pause_getI6242, pause_getI6249, pause_getI6257, pause_getI6266, pause_getI6274, pause_getI6278, pause_getI6286, pause_getI6291, pause_getI6295, pause_getI6300, pause_getI6306, pause_getI6312, pause_getI6319, pause_getI6326, pause_getI6337, pause_getI6341, pause_getI6346, pause_getI6353, pause_getI6360, pause_getI6369, pause_getI6373, pause_getI6385, pause_getI6393, pause_getI6397, pause_getI6401, pause_getI6409, pause_getI6414, pause_getI6418, pause_getI6429, pause_getI6433, pause_getI6437, pause_getI6446, pause_getI6454, pause_getI6458, pause_getI6466, pause_getI6471, pause_getI6475, pause_getI6479, pause_getI6489, pause_getI6497, pause_getI6501, pause_getI6509, pause_getI6514, pause_getI6518, pause_getI6522, pause_getI6532, pause_getI6540, pause_getI6544, pause_getI6552, pause_getI6557, pause_getI6561, pause_getI6566, pause_getI6585, pause_getI6596, pause_getI6601, pause_getI6610, pause_getI6618, pause_getI6622, pause_getI6630, pause_getI6635, pause_getI6639, pause_getI6643, pause_getI6653, pause_getI6661, pause_getI6665, pause_getI6673, pause_getI6678, pause_getI6682, pause_getI6686, pause_getI6695, pause_getI6703, pause_getI6707, pause_getI6715, pause_getI6720, pause_getI6724, pause_getI6729, pause_getI6748, pause_getI6758, pause_getI6762, pause_getI6771, pause_getI6779, pause_getI6783, pause_getI6791, pause_getI6796, pause_getI6800, pause_getI6804, pause_getI6814, pause_getI6822, pause_getI6826, pause_getI6834, pause_getI6839, pause_getI6843, pause_getI6847, pause_getI6856, pause_getI6864, pause_getI6868, pause_getI6876, pause_getI6881, pause_getI6885, pause_getI6890, pause_getI6909, pause_getI6919, pause_getI6923, pause_getI6933, pause_getI6941, pause_getI6945, pause_getI6953, pause_getI6958, pause_getI6962, pause_getI6972, pause_getI6976, pause_getI6987, pause_getI6991, pause_getII3379, pause_getII3398, pause_getII3405, pause_getII3419, pause_getII3426, pause_getII3434, pause_getII3444, pause_getII3451, pause_getII3460, pause_getII3472, pause_getII3479, pause_getII3488, pause_getII3495, pause_getII3506, pause_getII3512, pause_getII3520, pause_getII3529, pause_getII3537, pause_getII3541, pause_getII3549, pause_getII3554, pause_getII3558, pause_getII3569, pause_getII3573, pause_getII3582, pause_getII3588, pause_getII3598, pause_getII3606, pause_getII3610, pause_getII3618, pause_getII3623, pause_getII3627, pause_getII3639, pause_getII3645, pause_getII3657, pause_getII3669, pause_getII3676, pause_getII3685, pause_getII3691, pause_getII3696, pause_getII3707, pause_getII3713, pause_getII3726, pause_getII3734, pause_getII3738, pause_getII3742, pause_getII3750, pause_getII3755, pause_getII3759, pause_getII3763, pause_getII3771, pause_getII3779, pause_getII3783, pause_getII3791, pause_getII3796, pause_getII3800, pause_getII3811, pause_getII3815, pause_getII3826, pause_getII3830, pause_getII3841, pause_getII3845, pause_getII3854, pause_getII3862, pause_getII3866, pause_getII3870, pause_getII3878, pause_getII3883, pause_getII3887, pause_getII3898, pause_getII3902, pause_getII3913, pause_getII3917, pause_getII3926, pause_getII3934, pause_getII3938, pause_getII3942, pause_getII3950, pause_getII3955, pause_getII3959, pause_getII3970, pause_getII3974, pause_getII3985, pause_getII3989, pause_getII3998, pause_getII4006, pause_getII4010, pause_getII4014, pause_getII4022, pause_getII4027, pause_getII4031, pause_getII4035, pause_getII4044, pause_getII4052, pause_getII4056, pause_getII4064, pause_getII4069, pause_getII4073, pause_getII4077, pause_getII4082, pause_getII4095, pause_getII4099, pause_getII4110, pause_getII4118, pause_getII4122, pause_getII4126, pause_getII4134, pause_getII4139, pause_getII4143, pause_getII4157, pause_getII4161, pause_getII4170, pause_getII4178, pause_getII4182, pause_getII4186, pause_getII4194, pause_getII4199, pause_getII4203, pause_getII4208, pause_getII4221, pause_getII4225, pause_getII4234, pause_getII4242, pause_getII4246, pause_getII4250, pause_getII4258, pause_getII4263, pause_getII4267, pause_getII4272, pause_getII4285, pause_getII4289, pause_getII4298, pause_getII4306, pause_getII4310, pause_getII4314, pause_getII4322, pause_getII4327, pause_getII4331, pause_getII4336, pause_getII4349, pause_getII4353, pause_getII4362, pause_getII4370, pause_getII4374, pause_getII4378, pause_getII4386, pause_getII4391, pause_getII4395, pause_getII4405, pause_getII4412, pause_getII4427, pause_getII4431, pause_getII4442, pause_getII4446, pause_getII4455, pause_getII4463, pause_getII4467, pause_getII4471, pause_getII4479, pause_getII4484, pause_getII4488, pause_getII4498, pause_getII4505, pause_getII4520, pause_getII4524, pause_getII4535, pause_getII4539, pause_getII4548, pause_getII4556, pause_getII4560, pause_getII4564, pause_getII4572, pause_getII4577, pause_getII4581, pause_getII4591, pause_getII4598, pause_getII4613, pause_getII4617, pause_getII4628, pause_getII4632, pause_getII4643, pause_getII4651, pause_getII4655, pause_getII4659, pause_getII4667, pause_getII4672, pause_getII4676, pause_getII4715, pause_getII4722, pause_getII4739, pause_getII4743, pause_getII4754, pause_getII4758, pause_getII4767, pause_getII4775, pause_getII4779, pause_getII4783, pause_getII4791, pause_getII4796, pause_getII4800, pause_getII4819, pause_getII4823, pause_getII4834, pause_getII4838, pause_getII4847, pause_getII4855, pause_getII4859, pause_getII4863, pause_getII4871, pause_getII4876, pause_getII4880, pause_getII4898, pause_getII4902, pause_getII4913, pause_getII4917, pause_getII4926, pause_getII4934, pause_getII4938, pause_getII4942, pause_getII4950, pause_getII4955, pause_getII4959, pause_getII4977, pause_getII4981, pause_getII4992, pause_getII4996, pause_getII5005, pause_getII5013, pause_getII5017, pause_getII5021, pause_getII5029, pause_getII5034, pause_getII5038, pause_getII5056, pause_getII5060, pause_getII5071, pause_getII5075, pause_getII5084, pause_getII5092, pause_getII5096, pause_getII5100, pause_getII5108, pause_getII5113, pause_getII5117, pause_getII5135, pause_getII5139, pause_getII5150, pause_getII5154, pause_getII5163, pause_getII5171, pause_getII5175, pause_getII5179, pause_getII5187, pause_getII5192, pause_getII5196, pause_getII5205, pause_getII5213, pause_getII5217, pause_getII5221, pause_getII5229, pause_getII5234, pause_getII5238, pause_getII5252, pause_getII5256, pause_getII5264, pause_getII5272, pause_getII5279, pause_getII5286, pause_getII5291, pause_getII5300, pause_getII5306, pause_getII5311, pause_getII5315, pause_getII5327, pause_getII5333, pause_getII5344, pause_getII5351, pause_getII5360, pause_getII5367, pause_getII5377, pause_getII5384, pause_getII5401, pause_getII5405, pause_getII5417, pause_getII5423, pause_getII5432, pause_getII5440, pause_getII5444, pause_getII5448, pause_getII5456, pause_getII5461, pause_getII5465, pause_getII5471, pause_getII5478, pause_getII5485, pause_getII5490, pause_getII5506, pause_getII5512, pause_getII5521, pause_getII5529, pause_getII5533, pause_getII5537, pause_getII5545, pause_getII5550, pause_getII5554, pause_getII5566, pause_getII5572, pause_getII5602, pause_getII5606, pause_getII5614, pause_getII5620, pause_getII5641, pause_getII5645, pause_getII5653, pause_getII5658, pause_getII5662, pause_getII5666, pause_getII5670, pause_getII5678, pause_getII5683, pause_getII5687, pause_getII5699, pause_getII5705, pause_getII5716, pause_getII5723, pause_getII5732, pause_getII5738, pause_getII5750, pause_getII5756, pause_getII5767, pause_getII5774, pause_getII5783, pause_getII5789, pause_getII5801, pause_getII5807, pause_getII5818, pause_getII5825, pause_getII5834, pause_getII5840, pause_getII5852, pause_getII5858, pause_getII5868, pause_getII5875, pause_getII5884, pause_getII5890, pause_getII5894, pause_getII5904, pause_getII5912, pause_getII5916, pause_getII5924, pause_getII5929, pause_getII5933, pause_getII5937, pause_getII5949, pause_getII5956, pause_getII5962, pause_getII5972, pause_getII5979, pause_getII5987, pause_getII5996, pause_getII6004, pause_getII6008, pause_getII6016, pause_getII6021, pause_getII6025, pause_getII6030, pause_getII6036, pause_getII6047, pause_getII6051, pause_getII6061, pause_getII6068, pause_getII6076, pause_getII6085, pause_getII6093, pause_getII6097, pause_getII6105, pause_getII6110, pause_getII6114, pause_getII6119, pause_getII6125, pause_getII6133, pause_getII6137, pause_getII6147, pause_getII6155, pause_getII6159, pause_getII6167, pause_getII6172, pause_getII6176, pause_getII6180, pause_getII6189, pause_getII6197, pause_getII6201, pause_getII6209, pause_getII6214, pause_getII6218, pause_getII6229, pause_getII6233, pause_getII6243, pause_getII6250, pause_getII6258, pause_getII6267, pause_getII6275, pause_getII6279, pause_getII6287, pause_getII6292, pause_getII6296, pause_getII6301, pause_getII6307, pause_getII6313, pause_getII6320, pause_getII6327, pause_getII6338, pause_getII6342, pause_getII6347, pause_getII6354, pause_getII6361, pause_getII6370, pause_getII6374, pause_getII6386, pause_getII6394, pause_getII6398, pause_getII6402, pause_getII6410, pause_getII6415, pause_getII6419, pause_getII6430, pause_getII6434, pause_getII6438, pause_getII6447, pause_getII6455, pause_getII6459, pause_getII6467, pause_getII6472, pause_getII6476, pause_getII6480, pause_getII6490, pause_getII6498, pause_getII6502, pause_getII6510, pause_getII6515, pause_getII6519, pause_getII6523, pause_getII6533, pause_getII6541, pause_getII6545, pause_getII6553, pause_getII6558, pause_getII6562, pause_getII6567, pause_getII6586, pause_getII6597, pause_getII6602, pause_getII6611, pause_getII6619, pause_getII6623, pause_getII6631, pause_getII6636, pause_getII6640, pause_getII6644, pause_getII6654, pause_getII6662, pause_getII6666, pause_getII6674, pause_getII6679, pause_getII6683, pause_getII6687, pause_getII6696, pause_getII6704, pause_getII6708, pause_getII6716, pause_getII6721, pause_getII6725, pause_getII6730, pause_getII6749, pause_getII6759, pause_getII6763, pause_getII6772, pause_getII6780, pause_getII6784, pause_getII6792, pause_getII6797, pause_getII6801, pause_getII6805, pause_getII6815, pause_getII6823, pause_getII6827, pause_getII6835, pause_getII6840, pause_getII6844, pause_getII6848, pause_getII6857, pause_getII6865, pause_getII6869, pause_getII6877, pause_getII6882, pause_getII6886, pause_getII6891, pause_getII6910, pause_getII6920, pause_getII6924, pause_getII6934, pause_getII6942, pause_getII6946, pause_getII6954, pause_getII6959, pause_getII6963, pause_getII6973, pause_getII6977, pause_getII6988, pause_getII6992, pause_setI3370, pause_setI3384, pause_setI3392, pause_setI3413, pause_setI3438, pause_setI3466, pause_setI3524, pause_setI3532, pause_setI3544, pause_setI3561, pause_setI3593, pause_setI3601, pause_setI3613, pause_setI3630, pause_setI3648, pause_setI3663, pause_setI3721, pause_setI3729, pause_setI3745, pause_setI3766, pause_setI3774, pause_setI3786, pause_setI3803, pause_setI3818, pause_setI3833, pause_setI3849, pause_setI3857, pause_setI3873, pause_setI3890, pause_setI3905, pause_setI3921, pause_setI3929, pause_setI3945, pause_setI3962, pause_setI3977, pause_setI3993, pause_setI4001, pause_setI4017, pause_setI4039, pause_setI4047, pause_setI4059, pause_setI4087, pause_setI4105, pause_setI4113, pause_setI4129, pause_setI4149, pause_setI4165, pause_setI4173, pause_setI4189, pause_setI4213, pause_setI4229, pause_setI4237, pause_setI4253, pause_setI4277, pause_setI4293, pause_setI4301, pause_setI4317, pause_setI4341, pause_setI4357, pause_setI4365, pause_setI4381, pause_setI4399, pause_setI4419, pause_setI4434, pause_setI4450, pause_setI4458, pause_setI4474, pause_setI4492, pause_setI4512, pause_setI4527, pause_setI4543, pause_setI4551, pause_setI4567, pause_setI4585, pause_setI4605, pause_setI4620, pause_setI4638, pause_setI4646, pause_setI4662, pause_setI4731, pause_setI4746, pause_setI4762, pause_setI4770, pause_setI4786, pause_setI4811, pause_setI4826, pause_setI4842, pause_setI4850, pause_setI4866, pause_setI4890, pause_setI4905, pause_setI4921, pause_setI4929, pause_setI4945, pause_setI4969, pause_setI4984, pause_setI5000, pause_setI5008, pause_setI5024, pause_setI5048, pause_setI5063, pause_setI5079, pause_setI5087, pause_setI5103, pause_setI5127, pause_setI5142, pause_setI5158, pause_setI5166, pause_setI5182, pause_setI5200, pause_setI5208, pause_setI5224, pause_setI5244, pause_setI5318, pause_setI5338, pause_setI5371, pause_setI5393, pause_setI5408, pause_setI5427, pause_setI5435, pause_setI5451, pause_setI5497, pause_setI5516, pause_setI5524, pause_setI5540, pause_setI5557, pause_setI5575, pause_setI5594, pause_setI5623, pause_setI5629, pause_setI5636, pause_setI5648, pause_setI5673, pause_setI5690, pause_setI5710, pause_setI5741, pause_setI5761, pause_setI5792, pause_setI5812, pause_setI5843, pause_setI5862, pause_setI5899, pause_setI5907, pause_setI5919, pause_setI5940, pause_setI5966, pause_setI5991, pause_setI5999, pause_setI6011, pause_setI6039, pause_setI6055, pause_setI6080, pause_setI6088, pause_setI6100, pause_setI6142, pause_setI6150, pause_setI6162, pause_setI6184, pause_setI6192, pause_setI6204, pause_setI6221, pause_setI6237, pause_setI6262, pause_setI6270, pause_setI6282, pause_setI6333, pause_setI6365, pause_setI6381, pause_setI6389, pause_setI6405, pause_setI6425, pause_setI6442, pause_setI6450, pause_setI6462, pause_setI6485, pause_setI6493, pause_setI6505, pause_setI6528, pause_setI6536, pause_setI6548, pause_setI6606, pause_setI6614, pause_setI6626, pause_setI6649, pause_setI6657, pause_setI6669, pause_setI6691, pause_setI6699, pause_setI6711, pause_setI6767, pause_setI6775, pause_setI6787, pause_setI6810, pause_setI6818, pause_setI6830, pause_setI6852, pause_setI6860, pause_setI6872, pause_setI6929, pause_setI6937, pause_setI6949, pause_setI6968, pause_setI6983, pause_setI6995, pause_setI6999, pause_setI7003, pause_setI7007, pause_setI7011, pause_setI7015, pause_setII3371, pause_setII3385, pause_setII3393, pause_setII3414, pause_setII3439, pause_setII3467, pause_setII3525, pause_setII3533, pause_setII3545, pause_setII3562, pause_setII3594, pause_setII3602, pause_setII3614, pause_setII3631, pause_setII3649, pause_setII3664, pause_setII3722, pause_setII3730, pause_setII3746, pause_setII3767, pause_setII3775, pause_setII3787, pause_setII3804, pause_setII3819, pause_setII3834, pause_setII3850, pause_setII3858, pause_setII3874, pause_setII3891, pause_setII3906, pause_setII3922, pause_setII3930, pause_setII3946, pause_setII3963, pause_setII3978, pause_setII3994, pause_setII4002, pause_setII4018, pause_setII4040, pause_setII4048, pause_setII4060, pause_setII4088, pause_setII4106, pause_setII4114, pause_setII4130, pause_setII4150, pause_setII4166, pause_setII4174, pause_setII4190, pause_setII4214, pause_setII4230, pause_setII4238, pause_setII4254, pause_setII4278, pause_setII4294, pause_setII4302, pause_setII4318, pause_setII4342, pause_setII4358, pause_setII4366, pause_setII4382, pause_setII4400, pause_setII4420, pause_setII4435, pause_setII4451, pause_setII4459, pause_setII4475, pause_setII4493, pause_setII4513, pause_setII4528, pause_setII4544, pause_setII4552, pause_setII4568, pause_setII4586, pause_setII4606, pause_setII4621, pause_setII4639, pause_setII4647, pause_setII4663, pause_setII4732, pause_setII4747, pause_setII4763, pause_setII4771, pause_setII4787, pause_setII4812, pause_setII4827, pause_setII4843, pause_setII4851, pause_setII4867, pause_setII4891, pause_setII4906, pause_setII4922, pause_setII4930, pause_setII4946, pause_setII4970, pause_setII4985, pause_setII5001, pause_setII5009, pause_setII5025, pause_setII5049, pause_setII5064, pause_setII5080, pause_setII5088, pause_setII5104, pause_setII5128, pause_setII5143, pause_setII5159, pause_setII5167, pause_setII5183, pause_setII5201, pause_setII5209, pause_setII5225, pause_setII5245, pause_setII5319, pause_setII5339, pause_setII5372, pause_setII5394, pause_setII5409, pause_setII5428, pause_setII5436, pause_setII5452, pause_setII5498, pause_setII5517, pause_setII5525, pause_setII5541, pause_setII5558, pause_setII5576, pause_setII5595, pause_setII5624, pause_setII5630, pause_setII5637, pause_setII5649, pause_setII5674, pause_setII5691, pause_setII5711, pause_setII5742, pause_setII5762, pause_setII5793, pause_setII5813, pause_setII5844, pause_setII5863, pause_setII5900, pause_setII5908, pause_setII5920, pause_setII5941, pause_setII5967, pause_setII5992, pause_setII6000, pause_setII6012, pause_setII6040, pause_setII6056, pause_setII6081, pause_setII6089, pause_setII6101, pause_setII6143, pause_setII6151, pause_setII6163, pause_setII6185, pause_setII6193, pause_setII6205, pause_setII6222, pause_setII6238, pause_setII6263, pause_setII6271, pause_setII6283, pause_setII6334, pause_setII6366, pause_setII6382, pause_setII6390, pause_setII6406, pause_setII6426, pause_setII6443, pause_setII6451, pause_setII6463, pause_setII6486, pause_setII6494, pause_setII6506, pause_setII6529, pause_setII6537, pause_setII6549, pause_setII6607, pause_setII6615, pause_setII6627, pause_setII6650, pause_setII6658, pause_setII6670, pause_setII6692, pause_setII6700, pause_setII6712, pause_setII6768, pause_setII6776, pause_setII6788, pause_setII6811, pause_setII6819, pause_setII6831, pause_setII6853, pause_setII6861, pause_setII6873, pause_setII6930, pause_setII6938, pause_setII6950, pause_setII6969, pause_setII6984, pause_setII6996, pause_setII7000, pause_setII7004, pause_setII7008, pause_setII7012, pause_setII7016, q_wait3372, q_wait3380, q_wait3386, q_wait3394, q_wait3399, q_wait3406, q_wait3415, q_wait3420, q_wait3427, q_wait3435, q_wait3440, q_wait3445, q_wait3452, q_wait3461, q_wait3468, q_wait3473, q_wait3480, q_wait3489, q_wait3496, q_wait3507, q_wait3513, q_wait3521, q_wait3526, q_wait3530, q_wait3534, q_wait3538, q_wait3542, q_wait3546, q_wait3550, q_wait3555, q_wait3559, q_wait3563, q_wait3570, q_wait3574, q_wait3583, q_wait3589, q_wait3595, q_wait3599, q_wait3603, q_wait3607, q_wait3611, q_wait3615, q_wait3619, q_wait3624, q_wait3628, q_wait3632, q_wait3640, q_wait3646, q_wait3650, q_wait3658, q_wait3665, q_wait3670, q_wait3677, q_wait3686, q_wait3692, q_wait3697, q_wait3708, q_wait3714, q_wait3723, q_wait3727, q_wait3731, q_wait3735, q_wait3739, q_wait3743, q_wait3747, q_wait3751, q_wait3756, q_wait3760, q_wait3764, q_wait3768, q_wait3772, q_wait3776, q_wait3780, q_wait3784, q_wait3788, q_wait3792, q_wait3797, q_wait3801, q_wait3805, q_wait3812, q_wait3816, q_wait3820, q_wait3827, q_wait3831, q_wait3835, q_wait3842, q_wait3846, q_wait3851, q_wait3855, q_wait3859, q_wait3863, q_wait3867, q_wait3871, q_wait3875, q_wait3879, q_wait3884, q_wait3888, q_wait3892, q_wait3899, q_wait3903, q_wait3907, q_wait3914, q_wait3918, q_wait3923, q_wait3927, q_wait3931, q_wait3935, q_wait3939, q_wait3943, q_wait3947, q_wait3951, q_wait3956, q_wait3960, q_wait3964, q_wait3971, q_wait3975, q_wait3979, q_wait3986, q_wait3990, q_wait3995, q_wait3999, q_wait4003, q_wait4007, q_wait4011, q_wait4015, q_wait4019, q_wait4023, q_wait4028, q_wait4032, q_wait4036, q_wait4041, q_wait4045, q_wait4049, q_wait4053, q_wait4057, q_wait4061, q_wait4065, q_wait4070, q_wait4074, q_wait4078, q_wait4083, q_wait4089, q_wait4096, q_wait4100, q_wait4107, q_wait4111, q_wait4115, q_wait4119, q_wait4123, q_wait4127, q_wait4131, q_wait4135, q_wait4140, q_wait4144, q_wait4151, q_wait4158, q_wait4162, q_wait4167, q_wait4171, q_wait4175, q_wait4179, q_wait4183, q_wait4187, q_wait4191, q_wait4195, q_wait4200, q_wait4204, q_wait4209, q_wait4215, q_wait4222, q_wait4226, q_wait4231, q_wait4235, q_wait4239, q_wait4243, q_wait4247, q_wait4251, q_wait4255, q_wait4259, q_wait4264, q_wait4268, q_wait4273, q_wait4279, q_wait4286, q_wait4290, q_wait4295, q_wait4299, q_wait4303, q_wait4307, q_wait4311, q_wait4315, q_wait4319, q_wait4323, q_wait4328, q_wait4332, q_wait4337, q_wait4343, q_wait4350, q_wait4354, q_wait4359, q_wait4363, q_wait4367, q_wait4371, q_wait4375, q_wait4379, q_wait4383, q_wait4387, q_wait4392, q_wait4396, q_wait4401, q_wait4406, q_wait4413, q_wait4421, q_wait4428, q_wait4432, q_wait4436, q_wait4443, q_wait4447, q_wait4452, q_wait4456, q_wait4460, q_wait4464, q_wait4468, q_wait4472, q_wait4476, q_wait4480, q_wait4485, q_wait4489, q_wait4494, q_wait4499, q_wait4506, q_wait4514, q_wait4521, q_wait4525, q_wait4529, q_wait4536, q_wait4540, q_wait4545, q_wait4549, q_wait4553, q_wait4557, q_wait4561, q_wait4565, q_wait4569, q_wait4573, q_wait4578, q_wait4582, q_wait4587, q_wait4592, q_wait4599, q_wait4607, q_wait4614, q_wait4618, q_wait4622, q_wait4629, q_wait4633, q_wait4640, q_wait4644, q_wait4648, q_wait4652, q_wait4656, q_wait4660, q_wait4664, q_wait4668, q_wait4673, q_wait4677, q_wait4716, q_wait4723, q_wait4733, q_wait4740, q_wait4744, q_wait4748, q_wait4755, q_wait4759, q_wait4764, q_wait4768, q_wait4772, q_wait4776, q_wait4780, q_wait4784, q_wait4788, q_wait4792, q_wait4797, q_wait4801, q_wait4813, q_wait4820, q_wait4824, q_wait4828, q_wait4835, q_wait4839, q_wait4844, q_wait4848, q_wait4852, q_wait4856, q_wait4860, q_wait4864, q_wait4868, q_wait4872, q_wait4877, q_wait4881, q_wait4892, q_wait4899, q_wait4903, q_wait4907, q_wait4914, q_wait4918, q_wait4923, q_wait4927, q_wait4931, q_wait4935, q_wait4939, q_wait4943, q_wait4947, q_wait4951, q_wait4956, q_wait4960, q_wait4971, q_wait4978, q_wait4982, q_wait4986, q_wait4993, q_wait4997, q_wait5002, q_wait5006, q_wait5010, q_wait5014, q_wait5018, q_wait5022, q_wait5026, q_wait5030, q_wait5035, q_wait5039, q_wait5050, q_wait5057, q_wait5061, q_wait5065, q_wait5072, q_wait5076, q_wait5081, q_wait5085, q_wait5089, q_wait5093, q_wait5097, q_wait5101, q_wait5105, q_wait5109, q_wait5114, q_wait5118, q_wait5129, q_wait5136, q_wait5140, q_wait5144, q_wait5151, q_wait5155, q_wait5160, q_wait5164, q_wait5168, q_wait5172, q_wait5176, q_wait5180, q_wait5184, q_wait5188, q_wait5193, q_wait5197, q_wait5202, q_wait5206, q_wait5210, q_wait5214, q_wait5218, q_wait5222, q_wait5226, q_wait5230, q_wait5235, q_wait5239, q_wait5246, q_wait5253, q_wait5257, q_wait5265, q_wait5273, q_wait5280, q_wait5287, q_wait5292, q_wait5301, q_wait5307, q_wait5312, q_wait5316, q_wait5320, q_wait5328, q_wait5334, q_wait5340, q_wait5345, q_wait5352, q_wait5361, q_wait5368, q_wait5373, q_wait5378, q_wait5385, q_wait5395, q_wait5402, q_wait5406, q_wait5410, q_wait5418, q_wait5424, q_wait5429, q_wait5433, q_wait5437, q_wait5441, q_wait5445, q_wait5449, q_wait5453, q_wait5457, q_wait5462, q_wait5466, q_wait5472, q_wait5479, q_wait5486, q_wait5491, q_wait5499, q_wait5507, q_wait5513, q_wait5518, q_wait5522, q_wait5526, q_wait5530, q_wait5534, q_wait5538, q_wait5542, q_wait5546, q_wait5551, q_wait5555, q_wait5559, q_wait5567, q_wait5573, q_wait5577, q_wait5596, q_wait5603, q_wait5607, q_wait5615, q_wait5621, q_wait5625, q_wait5631, q_wait5638, q_wait5642, q_wait5646, q_wait5650, q_wait5654, q_wait5659, q_wait5663, q_wait5667, q_wait5671, q_wait5675, q_wait5679, q_wait5684, q_wait5688, q_wait5692, q_wait5700, q_wait5706, q_wait5712, q_wait5717, q_wait5724, q_wait5733, q_wait5739, q_wait5743, q_wait5751, q_wait5757, q_wait5763, q_wait5768, q_wait5775, q_wait5784, q_wait5790, q_wait5794, q_wait5802, q_wait5808, q_wait5814, q_wait5819, q_wait5826, q_wait5835, q_wait5841, q_wait5845, q_wait5853, q_wait5859, q_wait5864, q_wait5869, q_wait5876, q_wait5885, q_wait5891, q_wait5895, q_wait5901, q_wait5905, q_wait5909, q_wait5913, q_wait5917, q_wait5921, q_wait5925, q_wait5930, q_wait5934, q_wait5938, q_wait5942, q_wait5950, q_wait5957, q_wait5963, q_wait5968, q_wait5973, q_wait5980, q_wait5988, q_wait5993, q_wait5997, q_wait6001, q_wait6005, q_wait6009, q_wait6013, q_wait6017, q_wait6022, q_wait6026, q_wait6031, q_wait6037, q_wait6041, q_wait6048, q_wait6052, q_wait6057, q_wait6062, q_wait6069, q_wait6077, q_wait6082, q_wait6086, q_wait6090, q_wait6094, q_wait6098, q_wait6102, q_wait6106, q_wait6111, q_wait6115, q_wait6120, q_wait6126, q_wait6134, q_wait6138, q_wait6144, q_wait6148, q_wait6152, q_wait6156, q_wait6160, q_wait6164, q_wait6168, q_wait6173, q_wait6177, q_wait6181, q_wait6186, q_wait6190, q_wait6194, q_wait6198, q_wait6202, q_wait6206, q_wait6210, q_wait6215, q_wait6219, q_wait6223, q_wait6230, q_wait6234, q_wait6239, q_wait6244, q_wait6251, q_wait6259, q_wait6264, q_wait6268, q_wait6272, q_wait6276, q_wait6280, q_wait6284, q_wait6288, q_wait6293, q_wait6297, q_wait6302, q_wait6308, q_wait6314, q_wait6321, q_wait6328, q_wait6335, q_wait6339, q_wait6343, q_wait6348, q_wait6355, q_wait6362, q_wait6367, q_wait6371, q_wait6375, q_wait6383, q_wait6387, q_wait6391, q_wait6395, q_wait6399, q_wait6403, q_wait6407, q_wait6411, q_wait6416, q_wait6420, q_wait6427, q_wait6431, q_wait6435, q_wait6439, q_wait6444, q_wait6448, q_wait6452, q_wait6456, q_wait6460, q_wait6464, q_wait6468, q_wait6473, q_wait6477, q_wait6481, q_wait6487, q_wait6491, q_wait6495, q_wait6499, q_wait6503, q_wait6507, q_wait6511, q_wait6516, q_wait6520, q_wait6524, q_wait6530, q_wait6534, q_wait6538, q_wait6542, q_wait6546, q_wait6550, q_wait6554, q_wait6559, q_wait6563, q_wait6568, q_wait6587, q_wait6598, q_wait6603, q_wait6608, q_wait6612, q_wait6616, q_wait6620, q_wait6624, q_wait6628, q_wait6632, q_wait6637, q_wait6641, q_wait6645, q_wait6651, q_wait6655, q_wait6659, q_wait6663, q_wait6667, q_wait6671, q_wait6675, q_wait6680, q_wait6684, q_wait6688, q_wait6693, q_wait6697, q_wait6701, q_wait6705, q_wait6709, q_wait6713, q_wait6717, q_wait6722, q_wait6726, q_wait6731, q_wait6750, q_wait6760, q_wait6764, q_wait6769, q_wait6773, q_wait6777, q_wait6781, q_wait6785, q_wait6789, q_wait6793, q_wait6798, q_wait6802, q_wait6806, q_wait6812, q_wait6816, q_wait6820, q_wait6824, q_wait6828, q_wait6832, q_wait6836, q_wait6841, q_wait6845, q_wait6849, q_wait6854, q_wait6858, q_wait6862, q_wait6866, q_wait6870, q_wait6874, q_wait6878, q_wait6883, q_wait6887, q_wait6892, q_wait6911, q_wait6921, q_wait6925, q_wait6931, q_wait6935, q_wait6939, q_wait6943, q_wait6947, q_wait6951, q_wait6955, q_wait6960, q_wait6964, q_wait6970, q_wait6974, q_wait6978, q_wait6985, q_wait6989, q_wait6993, q_wait6997, q_wait7001, q_wait7005, q_wait7009, q_wait7013, q_wait7017);
  signal state_var7021: t_state_var7021;
  type array_value_32 is array (natural range <>) of value(0 to 31);
  type array_value_108 is array (natural range <>) of value(0 to 107);
  signal \$10695_limit\ : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$$10695_limit_value\ : value(0 to 31);
  signal \$$10695_limit_ptr\ : natural range 0 to 0;
  signal \$$10695_limit_ptr_write\ : natural range 0 to 0;
  signal \$$10695_limit_write\ : value(0 to 31);
  signal \$$10695_limit_write_request\ : std_logic := '0';
  signal \$10696_ram\ : array_value_108(0 to 9999) := (others => (others => '0'));
  signal \$$10696_ram_value\ : value(0 to 107);
  signal \$$10696_ram_ptr\ : natural range 0 to 9999;
  signal \$$10696_ram_ptr_write\ : natural range 0 to 9999;
  signal \$$10696_ram_write\ : value(0 to 107);
  signal \$$10696_ram_write_request\ : std_logic := '0';
  signal \$10697_stack\ : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$$10697_stack_value\ : value(0 to 31);
  signal \$$10697_stack_ptr\ : natural range 0 to 0;
  signal \$$10697_stack_ptr_write\ : natural range 0 to 0;
  signal \$$10697_stack_write\ : value(0 to 31);
  signal \$$10697_stack_write_request\ : std_logic := '0';
  signal \$10698_heap\ : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$$10698_heap_value\ : value(0 to 31);
  signal \$$10698_heap_ptr\ : natural range 0 to 0;
  signal \$$10698_heap_ptr_write\ : natural range 0 to 0;
  signal \$$10698_heap_write\ : value(0 to 31);
  signal \$$10698_heap_write_request\ : std_logic := '0';
  signal \$10699_symtbl\ : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$$10699_symtbl_value\ : value(0 to 31);
  signal \$$10699_symtbl_ptr\ : natural range 0 to 0;
  signal \$$10699_symtbl_ptr_write\ : natural range 0 to 0;
  signal \$$10699_symtbl_write\ : value(0 to 31);
  signal \$$10699_symtbl_write_request\ : std_logic := '0';
  signal \$10700_pc\ : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$$10700_pc_value\ : value(0 to 31);
  signal \$$10700_pc_ptr\ : natural range 0 to 0;
  signal \$$10700_pc_ptr_write\ : natural range 0 to 0;
  signal \$$10700_pc_write\ : value(0 to 31);
  signal \$$10700_pc_write_request\ : std_logic := '0';
  signal \$10701_pos\ : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$$10701_pos_value\ : value(0 to 31);
  signal \$$10701_pos_ptr\ : natural range 0 to 0;
  signal \$$10701_pos_ptr_write\ : natural range 0 to 0;
  signal \$$10701_pos_write\ : value(0 to 31);
  signal \$$10701_pos_write_request\ : std_logic := '0';
  signal \$10702_brk\ : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$$10702_brk_value\ : value(0 to 31);
  signal \$$10702_brk_ptr\ : natural range 0 to 0;
  signal \$$10702_brk_ptr_write\ : natural range 0 to 0;
  signal \$$10702_brk_write\ : value(0 to 31);
  signal \$$10702_brk_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$$10695_limit_write_request\ = '1' then
                    \$10695_limit\(\$$10695_limit_ptr_write\) <= \$$10695_limit_write\;
                  else
                   \$$10695_limit_value\ <= \$10695_limit\(\$$10695_limit_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$$10696_ram_write_request\ = '1' then
                    \$10696_ram\(\$$10696_ram_ptr_write\) <= \$$10696_ram_write\;
                  else
                   \$$10696_ram_value\ <= \$10696_ram\(\$$10696_ram_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$$10697_stack_write_request\ = '1' then
                    \$10697_stack\(\$$10697_stack_ptr_write\) <= \$$10697_stack_write\;
                  else
                   \$$10697_stack_value\ <= \$10697_stack\(\$$10697_stack_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$$10698_heap_write_request\ = '1' then
                    \$10698_heap\(\$$10698_heap_ptr_write\) <= \$$10698_heap_write\;
                  else
                   \$$10698_heap_value\ <= \$10698_heap\(\$$10698_heap_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$$10699_symtbl_write_request\ = '1' then
                    \$10699_symtbl\(\$$10699_symtbl_ptr_write\) <= \$$10699_symtbl_write\;
                  else
                   \$$10699_symtbl_value\ <= \$10699_symtbl\(\$$10699_symtbl_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$$10700_pc_write_request\ = '1' then
                    \$10700_pc\(\$$10700_pc_ptr_write\) <= \$$10700_pc_write\;
                  else
                   \$$10700_pc_value\ <= \$10700_pc\(\$$10700_pc_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$$10701_pos_write_request\ = '1' then
                    \$10701_pos\(\$$10701_pos_ptr_write\) <= \$$10701_pos_write\;
                  else
                   \$$10701_pos_value\ <= \$10701_pos\(\$$10701_pos_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$$10702_brk_write_request\ = '1' then
                    \$10702_brk\(\$$10702_brk_ptr_write\) <= \$$10702_brk_write\;
                  else
                   \$$10702_brk_value\ <= \$10702_brk\(\$$10702_brk_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable result3362 : value(0 to 1) := (others => '0');
      variable \$13500_list_tail2653266_result\, \$v5330\, \$v3502\, 
               \$11663\, \$v4508\, \$v6357\, \$v6226\, \$v4439\, \$12777_x\, 
               \$v5746\, \$v6903\, \$v6064\, \$15076_new_rib\, \$v6745\, 
               \$v5984\, \$v5728\, \$v4706\, \$14542_new_rib\, \$v5797\, 
               \$11437_loop3073170_result\, \$v4989\, \$11911\, \$v3895\, 
               \$v5474\, \$v5242\, \$v5887\, \$11556_z\, \$10839_s\, 
               \$v4831\, \$v5871\, \$12428_y\, \$11219\, \$12877_x\, 
               \$12686_y\, \$13666\, \$v5848\, \$v5880\, \$v5562\, \$v3703\, 
               \$v5982\, \$11223\, \$v5495\, \$v5387\, \$v5569\, \$v3491\, 
               \$v6756\, \$v3808\, \$v3484\, \$v4085\, \$15475_end_rib\, 
               \$v3672\, \$v5821\, \$v3585\, \$v5391\, \$v5356\, \$11809\, 
               \$14840\, \$v5502\, \$11548_y\, \$v3447\, \$v4718\, \$v6073\, 
               \$v3578\, \$v4751\, \$11736_x\, \$v4681\, \$15467_str_rib\, 
               \$v5726\, \$v4532\, \$v5260\, \$v5975\, \$v4339\, \$v5830\, 
               \$13085_y\, \$v5275\, \$10828_c2_rib\, \$12305_y\, \$v5068\, 
               \$v4709\, \$v6033\, \$v5837\, \$12678_x\, \$12543_x\, 
               \$14648_ty\, \$v3463\, \$v6122\, \$v4346\, \$15303_str_rib\, 
               \$v5959\, \$v4424\, \$v5053\, \$12785_y\, \$v6579\, \$v4147\, 
               \$12420_x\, \$15068_opnd\, \$12985_y\, \$10897_k\, \$v5294\, 
               \$v5147\, \$v4701\, \$v5354\, \$v3422\, 
               \$14863_list_tail2653331_result\, \$v6255\, \$v5125\, 
               \$v4415\, \$11328_cont\, \$v6246\, \$v4729\, \$12105\, 
               \$v4967\, \$v3375\, \$v3660\, \$13295\, \$v3456\, \$v3653\, 
               \$13596_v\, \$v5380\, \$v6304\, \$v4601\, \$v4691\, \$v3429\, 
               \$v4888\, \$v5481\, \$v5702\, \$v5413\, \$v3910\, \$13222\, 
               \$13405\, \$v5828\, \$v4727\, \$12786\, \$v4218\, \$v5363\, 
               \$v3681\, \$12297_x\, \$v5509\, \$11814\, \$v5323\, \$v6575\, 
               \$v3431\, \$v3475\, \$14533_opnd\, \$v6570\, \$13086\, 
               \$v4625\, \$v3838\, \$v4154\, \$v4092\, \$v5779\, \$v5786\, 
               \$v4275\, \$12182_y\, \$13077_x\, 
               \$13318_list_tail2653256_result\, \$v5267\, \$v5804\, 
               \$12977_x\, \$14656_proc_rib\, \$v4517\, \$13221\, \$v5719\, 
               \$12687\, \$v4686\, \$v6316\, \$v5493\, \$v3454\, 
               \$14652_code_proc_rib\, \$v3498\, \$v4974\, \$13813\, 
               \$v3401\, \$v3688\, \$v4816\, \$v6582\, \$v4910\, \$v5617\, 
               \$13689_list_tail2653276_result\, \$v5770\, \$v5695\, 
               \$v3566\, \$10738_main_rib\, \$v5585\, \$v5303\, \$v3679\, 
               \$12986\, \$v4809\, \$v5389\, \$v3982\, \$v5296\, \$v6253\, 
               \$12551_y\, \$11036_loop3073149_result\, \$11967\, \$v3710\, 
               \$v4501\, \$v4510\, \$v5347\, \$15642_end_rib\, \$v4689\, 
               \$v6752\, \$v5753\, \$v6917\, \$v5855\, 
               \$14996_list_tail2653334_result\, \$v6589\, \$v4736\, 
               \$v3482\, \$v3517\, \$12174_x\, \$v5249\, \$v3389\, \$v6899\, 
               \$v4594\, \$15634_str_rib\, \$v3509\, \$v3823\, \$v6742\, 
               \$13174\, \$v3642\, \$14973\, \$v4282\, \$v5599\, \$v4807\, 
               \$12886\, \$11540_x\, \$v3410\, \$v4886\, \$v6044\, \$v5398\, 
               \$v4408\, \$v4696\, \$v3408\, \$v5044\, \$v6350\, \$v5878\, 
               \$v4965\, \$10818_proc\, \$v6738\, \$v5589\, \$v5580\, 
               \$v4895\, \$v6906\, \$v6913\, \$v5132\, 
               \$11196_loop2913158_result\, \$12885_y\, \$v5123\, \$v4699\, 
               \$v3635\, \$15267\, \$v6593\, \$12036\, \$v5420\, \$v5046\, 
               \$15311_end_rib\, \$14667_new_rib\, \$v6733\, \$v5735\, 
               \$v4711\, \$v6323\, \$v4417\, \$v3967\, \$v3699\, \$v5777\, 
               \$13446\, \$v5610\, \$v6894\, \$v4603\, \$v5952\, \$v3382\, 
               \$v4725\, \$v5945\, \$v5592\, \$11564_r\, \$v5282\, \$v4610\, 
               \$v3718\, \$v6071\, \$v4211\, \$v6130\ : value(0 to 35) := (others => '0');
      variable \$14939_get_int268_arg\, \$15788_get_int268_arg\, 
               \$14897_get_int268_arg\ : value(0 to 32) := (others => '0');
      variable \$11437_loop3073170_arg\, \$11036_loop3073149_arg\ : value(0 to 36) := (others => '0');
      variable \$14511_loop311_arg\ : value(0 to 102) := (others => '0');
      variable \$15555_len_aux3143354_arg\, \$13318_list_tail2653256_arg\, 
               \$14863_list_tail2653331_arg\, \$14996_list_tail2653334_arg\, 
               \$15724_len_aux3143361_arg\, \$13500_list_tail2653266_arg\, 
               \$13689_list_tail2653276_arg\, \$15391_len_aux3143348_arg\ : value(0 to 68) := (others => '0');
      variable \$v3432\, \$v5946\, \$v6317\, \$v5590\, \$v5399\, \$v4808\, 
               \$v5729\, \$v5787\, \$v5798\, \$v3476\, \$v4212\, \$v3409\, 
               \$v4283\, \$v6074\, \$v5581\, \$v5381\, \$v3983\, \$v5297\, 
               \$v6576\, \$v5805\, \$v3510\, \$v6123\, \$v5268\, \$v6571\, 
               \$v4737\, \$v6904\, \$v4626\, \$v5510\, \$v3643\, \$v5829\, 
               \$v4889\, \$v3455\, \$v5045\, \$v5475\, \$v5881\, \$v5126\, 
               \$v5983\, \$v3636\, \$v3457\, \$v5421\, \$v5720\, \$v6045\, 
               \$v6580\, \$v4810\, \$v4702\, \$v6305\, \$v5276\, \$v4990\, 
               \$v6072\, \$v4911\, \$v5976\, \$v4347\, \$v5133\, \$v4602\, 
               \$v5727\, \$v4155\, \$v5563\, \$v5822\, \$v3567\, \$v5696\, 
               \$v3376\, \$v4502\, \$v4712\, \$v5872\, \$v3896\, \$v3661\, 
               \$v4086\, \$v6918\, \$v3448\, \$v5482\, \$v5390\, \$v3689\, 
               \$v5747\, \$v6590\, \$v5780\, \$v5047\, \$v3430\, \$v5570\, 
               \$v3383\, \$v5618\, \$v5496\, \$v5778\, \$v4726\, \$v5324\, 
               \$v3499\, \$v5856\, \$v6254\, \$v5771\, \$v5124\, \$v5392\, 
               \$v6739\, \$v4817\, \$v4595\, \$v5831\, \$v3483\, \$v5388\, 
               \$v3503\, \$v5348\, \$v5331\, \$v5261\, \$v3682\, \$v3411\, 
               \$v4728\, \$v4611\, \$v6351\, \$v5586\, \$v3719\, \$v4511\, 
               \$v4340\, \$v5953\, \$v4509\, \$v4966\, \$v4687\, \$v5754\, 
               \$v4896\, \$v5503\, \$v6757\, \$v4093\, \$v5600\, \$v5355\, 
               \$v5879\, \$v3680\, \$v4968\, \$v4697\, \$v3704\, \$v3911\, 
               \$v3586\, \$v5593\, \$v6895\, \$v3700\, \$v4707\, \$v4219\, 
               \$v4752\, \$v5736\, \$v4730\, \$v5283\, \$v5888\, \$v6358\, 
               \$v3485\, \$v5960\, \$v6583\, \$v4533\, \$v6324\, \$v3423\, 
               \$v5849\, \$v5243\, \$v5494\, \$v4719\, \$v6907\, \$v4690\, 
               \$v6227\, \$v3711\, \$v6247\, \$v5304\, \$v4832\, \$v6256\, 
               \$v3464\, \$v3518\, \$v6734\, \$v4700\, \$v3654\, \$v4887\, 
               \$v5295\, \$v4440\, \$v5054\, \$v6743\, \$v6900\, \$v4418\, 
               \$v4682\, \$v3968\, \$v6594\, \$v3579\, \$v4518\, \$v3492\, 
               \$v3673\, \$v6065\, \$v6034\, \$v3839\, \$v5611\, \$v6753\, 
               \$v5357\, \$v4975\, \$v5985\, \$v5148\, \$v4409\, \$v4425\, 
               \$v3390\, \$v5069\, \$v6914\, \$v6131\, \$v6746\, \$v4148\, 
               \$v3809\, \$v5250\, \$v4276\, \$v5838\, \$v5364\, \$v4692\, 
               \$v4416\, \$v5703\, \$v5414\, \$v3402\, \$v3824\, \$v4710\, 
               \$v4604\ : value(0 to 3) := (others => '0');
      variable \$11196_loop2913158_arg\ : value(0 to 72) := (others => '0');
      variable \$15240_loop23133355_arg\ : value(0 to 41) := (others => '0');
      variable \$15217_loop1312_arg\ : value(0 to 37) := (others => '0');
      variable \$v3428\, \$v5547\, rdy3366, \$v5535\, \$v3864\, \$v6932\, 
               \$v4869\, \$v6063\, \$v4397\, \$v6944\, \$v6867\, \$v5215\, 
               \$v6488\, \$v3868\, \$v5914\, \$v5886\, \$v6310\, \$v5854\, 
               \$v4829\, \$v5668\, \$v6879\, \$v3828\, \$v6145\, \$v6465\, 
               \$v4008\, \$v3817\, \$v5902\, \$v4296\, \$v5910\, \$v5681\, 
               \$v4012\, \$v6634\, \$v4477\, \$v4444\, \$v4575\, \$v5680\, 
               \$v5877\, \$v6952\, \$v5660\, \$v7002\, \$v5676\, \$v4261\, 
               \$v5672\, \$v6564\, \$v6975\, \$v6191\, \$v3952\, \$v4717\, 
               \$v5236\, \$v4657\, \$v5115\, \$v6915\, \$v6412\, \$v5219\, 
               \$v6966\, \$14511_loop311_result\, \$v5758\, \$v5939\, 
               \$15217_loop1312_result\, \$v5906\, \$v4269\, \$v5718\, 
               \$v6153\, \$v5062\, \$v4789\, \$v6170\, \$v5106\, \$11912\, 
               \$v6157\, \$12552\, \$v3497\, \$v6032\, \$v4987\, \$v5473\, 
               \$v5403\, \$v3647\, \$v6807\, \$v4024\, \$v6290\, \$v6833\, 
               \$v4526\, \$v5110\, \$v5713\, \$v4108\, \$v5500\, \$v4583\, 
               \$v3709\, \$v5803\, \$v5989\, \$v5483\, \$v3659\, \$v4600\, 
               \$v5531\, \$v5922\, \$v5701\, \$v4372\, \$v6422\, \$v6672\, 
               \$v4256\, \$v5111\, \$v6231\, \$v6368\, \$v5341\, \$v4137\, 
               \$v4670\, \$v6377\, \$v6457\, \$v4630\, \$v5274\, \$v5190\, 
               \$v3744\, \$v3852\, \$v6638\, \$v4665\, \$v6212\, \$v5827\, 
               \$v6315\, \$v6735\, \$v3972\, \$v5791\, \$v3813\, \$v6332\, 
               \$15563\, \$v6604\, \$v4857\, \$v5556\, \$v6187\, \$v6990\, 
               \$v3724\, \$v5051\, \$v5353\, \$v4953\, \$v5396\, \$v4216\, 
               \$v4836\, \$11448\, \$v3732\, \$v6099\, \$v6285\, \$15564\, 
               \$v5454\, \$v5156\, \$v3400\, \$v4983\, \$v5548\, \$v4128\, 
               \$v4794\, \$v4550\, \$v4608\, \$v3469\, \$v5231\, \$v4422\, 
               \$v6754\, \$v4252\, \$v6685\, \$v7014\, \$v3924\, \$v4168\, 
               \$v4016\, \$v6135\, \$v3716\, \$11047\, \$v4000\, \$v6689\, 
               \$v6216\, \$v6859\, \$v3552\, \$v5102\, \$v5597\, \$v5508\, 
               \$v6875\, \$v4932\, \$v5560\, \$v6795\, \$v4457\, \$v4388\, 
               \$v5335\, \$v7010\, \$v6359\, \$v3940\, \$v5141\, \$v4558\, 
               \$v4825\, \$v6449\, \$v4994\, \$v6325\, \$v6714\, \$v6893\, 
               \$v3793\, \$v4025\, \$v3769\, \$v5734\, rdy3363, \$v4465\, 
               \$v4101\, \$v5725\, \$v3527\, \$v5463\, \$v3843\, \$v5492\, 
               \$v3531\, \$v3753\, \$v6521\, \$v5073\, \$v4141\, \$v3773\, 
               \$v4172\, \$v5198\, \$v3715\, \$v6718\, \$v4861\, \$v3736\, 
               \$v6922\, \$v6660\, \$v6535\, \$v5552\, \$v4802\, \$v6940\, 
               \$v5040\, \$v6965\, \$v4957\, \$v3381\, \$v3928\, \$v4380\, 
               \$v5365\, \$v6646\, \$v4360\, \$v4678\, \$v4260\, \$v4653\, 
               \$v6863\, \$v6846\, \$v4042\, \$v4915\, \$v4546\, \$v5011\, 
               \$v6245\, \$v3678\, \$v5036\, \$v6525\, \$v4554\, \$v6421\, 
               \$v6424\, \$v6994\, \$v6799\, \$v6817\, \$v6912\, \$v5077\, 
               \$v6289\, \$v3373\, \$v5098\, \$v3535\, \$v4180\, \$v5523\, 
               \$v3701\, \$14481_decode_loop310_result\, \$v3543\, \$v5090\, 
               \$v6979\, \$v5169\, \$v6998\, \$v6961\, \$v6478\, \$v6388\, 
               \$v6400\, \$v4402\, \$v6569\, \$v4090\, \$v3387\, \$v5809\, 
               \$v5189\, \$v5266\, \$15240_loop23133355_result\, \$v3915\, 
               \$v4777\, \$v6116\, \$v5007\, \$v3980\, \$v4495\, \$v3860\, 
               \$v6364\, \$v6782\, \$v3490\, \$v6182\, \$v6165\, \$v6252\, 
               \$v5568\, \$v4669\, \$v6269\, \$v4724\, \$v4570\, \$15733\, 
               \$v6794\, \$v5329\, \$v4645\, \$v4944\, \$v6112\, \$v3500\, 
               \$v6609\, \$v6681\, \$12597\, \$v3752\, \$v5346\, \$v4473\, 
               \$v3514\, \$v3551\, \$v5317\, \$v6825\, \$v4355\, \$v3836\, 
               \$v3600\, \$v6445\, \$v4308\, \$v4588\, \$v4210\, \$v4364\, 
               \$v6203\, \$v6803\, \$v3539\, \$v5130\, \$v5173\, \$v3893\, 
               \$v6706\, \$12598\, \$v6303\, \$v4469\, \$v3991\, \$v3416\, 
               \$v5223\, \$v6555\, \$v3621\, \$v6710\, \$v4623\, \$v5943\, 
               \$v7018\, \$v6413\, \$v4197\, \$v6492\, \$v6676\, \$v4878\, 
               \$v4236\, \$v6392\, \$v5321\, \$v6108\, \$v6621\, \$v6838\, 
               \$v5308\, \$v6161\, \$v4745\, result3365, \$v6668\, \$v4908\, 
               \$v6235\, \$v6633\, \$v3633\, \$v6664\, \$v5288\, \$v6298\, 
               \$v4579\, \$v4936\, \$v6936\, \$v5058\, \$v3547\, \$v3965\, 
               \$v4845\, \$v4287\, \$v6560\, \$v4481\, \$v4205\, \$v3596\, 
               \$v6091\, \$v5764\, \$v6273\, \$v4265\, \$v4853\, \$v6372\, 
               \$v6652\, \$v5119\, \$v6376\, \$v6572\, \$v4979\, \$v5632\, 
               \$v4058\, \$v4769\, \$v6404\, \$v3748\, \$v4033\, \$v6469\, 
               \$v5776\, \$v6309\, \$v4900\, \$v6336\, \$v3889\, \$v4329\, 
               \$v6625\, \$v3932\, \$v5892\, \$v6384\, \$v6139\, \$v4515\, 
               \$v6019\, \$v4046\, \$v6821\, \$v4037\, \$v3953\, \$v5643\, 
               \$v4961\, \$v4020\, \$v6127\, \$v4693\, \$v3900\, \$v6408\, 
               \$v3395\, \$v6957\, \$v3936\, \$v5896\, \$v6349\, \$v4244\, 
               \$v5438\, \$v6224\, \$v6010\, \$v3687\, \$v5981\, \$v6396\, 
               \$v3806\, \$v4840\, \$v4291\, \$v6613\, \$v6107\, \$v5240\, 
               \$v4566\, \$v4152\, \$v5480\, \$v5207\, \$v6432\, \$v3872\, 
               \$v5165\, \$v4919\, \$v3740\, \$v6888\, \$v6018\, \$v4522\, 
               \$v5258\, \$v5527\, \$v5842\, \$v6871\, \$15400\, \$v3880\, 
               \$v3728\, \$v5926\, \$v6837\, \$v4145\, \$v5974\, \$v6006\, 
               \$v7006\, \$v3765\, \$v5740\, \$v6770\, \$v6727\, \$v3620\, 
               \$v6850\, \$v6539\, \$v6281\, \$v6169\, \$v6331\, \$v3560\, 
               \$v6195\, \$v5969\, \$v6556\, \$v3976\, \$v6842\, \$v3885\, 
               \$v5820\, \$v4223\, \$v6698\, \$v4316\, \$v4649\, \$v4765\, 
               \$v4304\, \$v6260\, \$v4344\, \$v4785\, \$v3608\, \$15732\, 
               \$v3856\, \$v5927\, \$v5302\, \$v4124\, \$v6220\, \$v4849\, 
               \$v6363\, \$v5374\, \$v3948\, \$v5918\, \$v3832\, \$v6440\, 
               \$v5177\, \$v6178\, \$v3789\, \$v3436\, \$v6517\, \$v3944\, 
               \$v6417\, \$v6926\, \$15399\, \$v5211\, \$v6083\, \$v5362\, 
               \$v5578\, \$v3908\, \$v6774\, \$v5626\, \$v6423\, \$v4232\, 
               \$v6174\, \$v3446\, \$v4333\, \$v3757\, \$v4448\, \$v4530\, 
               \$v5032\, \$v6778\, \$v6294\, \$v5181\, \$v5459\, \$v5685\, 
               \$v3575\, \$v3441\, \$v3693\, \$v3522\, \$v6340\, \$v4066\, 
               \$v6948\, \$v5785\, \$v4461\, \$v5543\, \$v6002\, \$v6982\, 
               \$v6322\, \$v4312\, \$v5094\, \$v6813\, \$v4075\, \$v3584\, 
               \$v4320\, \$v4227\, \$v4240\, \$v6677\, \$v6149\, \$v5689\, 
               \$v6504\, \$v3481\, \$v6531\, \$v3556\, \$v5185\, \$v5293\, 
               \$v6436\, \$v3671\, \$v5313\, \$v5023\, \$13814\, \$v4192\, 
               \$v4507\, \$v5434\, \$v4482\, \$v5411\, \$v5194\, \$v3616\, 
               \$v6378\, \$v5744\, \$v3612\, \$v3515\, \$v4873\, \$v6956\, 
               \$10778_run286_result\, \$v3576\, \$v3881\, \$v5865\, 
               \$v6474\, \$v4948\, \$v3564\, \$v4274\, \$v6617\, \$v5693\, 
               \$v6981\, \$v4773\, \$v5145\, \$v4132\, \$v4562\, \$v5998\, 
               \$v6719\, \$v3590\, \$v3421\, \$v6053\, \$v5707\, \$v6588\, 
               \$v5254\, \$v4972\, \$v5622\, \$v4793\, \$v5386\, \$v5964\, 
               \$v3781\, \$v6829\, \$v6880\, \$v5664\, \$v4821\, \$v6356\, 
               \$v6694\, \$v4940\, \$v5425\, \$v6329\, \$v5066\, \$v6790\, 
               \$v5309\, \$v6023\, \$v4615\, \$v4882\, \$v6087\, \$v5446\, 
               \$v6547\, \$v4376\, \$v3651\, \$v5487\, \$v4196\, \$v6786\, 
               \$v7020\, \$v4324\, \$v3821\, \$v4865\, \$v4593\, \$v5086\, 
               \$v6543\, \$v6765\, \$v3761\, \$v5227\, \$v5082\, \$v6042\, 
               \$v4429\, \$v4062\, \$v5015\, \$v5574\, \$v5281\, \$v6049\, 
               \$v5994\, \$v3785\, \$v4998\, \$v3802\, \$v4338\, \$v4071\, 
               \$v5608\, \$v6265\, \$v4389\, \$v4201\, \$v5419\, \$v5769\, 
               \$v6971\, \$v6207\, \$v5467\, \$v3794\, \$v3625\, \$v6121\, 
               \$v3666\, \$v4176\, \$v3474\, \$v5003\, \$v4407\, \$v6014\, 
               \$v6656\, \$11323\, \$v5656\, \$v3777\, \$v4537\, \$v6761\, 
               \$v4619\, \$v3961\, \$v4163\, \$v4159\, \$v4490\, \$v6629\, 
               \$v4500\, \$v5379\, \$v3407\, \$v6103\, \$v6453\, \$v4384\, 
               \$v5651\, \$v6751\, \$v6482\, \$v3996\, \$v4112\, \$v5450\, 
               \$v5161\, \$v4188\, \$v5031\, \$v4924\, \$v4893\, \$v4067\, 
               \$v4184\, \$v4368\, \$v5647\, \$v6896\, \$v6344\, \$v4541\, 
               \$v4453\, \$v5795\, \$v4756\, \$v6277\, \$v4248\, \$v6702\, 
               \$v6986\, \$v3987\, \$v5846\, \$v4798\, \$v5815\, \$v5951\, 
               \$v6428\, \$v5203\, \$v4661\, \$v4574\, \$v6461\, \$v5870\, 
               \$v6884\, \$v5539\, \$v3641\, \$v4414\, \$v5860\, \$10840\, 
               \$v5027\, \$v5247\, \$v3904\, \$v5519\, \$v5284\, \$v4928\, 
               \$v3698\, \$v6551\, \$v4433\, \$v4393\, \$v4641\, \$v6038\, 
               \$v4097\, \$v6723\, \$v4634\, \$v5514\, \$v6513\, \$v3629\, 
               \$v5430\, \$v5958\, \$v3604\, \$v4674\, \$v6058\, \$v3876\, 
               \$v5639\, \$v3957\, \$v3847\, \$v6732\, \$v4280\, \$v4116\, 
               \$v4136\, \$v6211\, \$v5582\, \$v6095\, \$v6591\, \$v6508\, 
               \$v5604\, \$v4351\, \$v5655\, \$v4734\, \$v4054\, \$v4004\, 
               \$v3508\, \$v6599\, \$v4029\, \$v4952\, \$v6470\, \$v6496\, 
               \$v6500\, \$v6078\, \$v6027\, \$v4300\, \$v6967\, \$v5019\, 
               \$v3919\, \$v3798\, \$v3453\, \$v5931\, \$v5137\, \$v5935\, 
               \$v5836\, \$v6855\, \$v5407\, \$v4084\, \$v5752\, \$v4050\, 
               \$v4437\, \$14659\, \$v4741\, \$v5369\, \$v3462\, \$v4486\, 
               \$v4749\, \$v4760\, \$v6199\, \$v6128\, \$v4904\, \$v5616\, 
               \$v6240\, \$v4781\, \$v5458\, \$v4814\, \$v4703\, \$v5152\, 
               \$v4120\, \$v4874\, \$v4079\, \$v6070\, \$v6512\, \$v4325\, 
               \$v5442\, \$v5232\, \$v3571\, \$v6642\ : value(0 to 0) := (others => '0');
      variable \$14682\, \$11443\, \$13547\, \$12872\, \$11100\, \$11804\, 
               \$13327\, \$11535\, \$11048\, \$11380\, \$12226\, \$11709\, 
               \$15734\, \$13216\, \$11149\, \$10848\, \$13460\, \$11551\, 
               \$14872\, \$13967\, \$11543\, \$14301\, \$10750\, \$12415\, 
               \$14683\, \$12587\, \$13296\, \$12972\, \$11658\, \$12980\, 
               \$12169\, \$14662\, \$10721\, \$15091\, \$10900\, \$13832\, 
               \$14080\, \$11962\, \$10814\, \$12473\, \$14643\, \$13509\, 
               \$12300\, \$13750\, \$10726\, \$14558\, \$10981\, \$12031\, 
               \$14974\, \$11333\, \$15755\, \$10793\, \$10980\, \$12880\, 
               \$11214\, \$13461\, \$15071\, \$13667\, \$14017\, \$11449\, 
               \$13546\, \$11148\, \$13607\, \$11042\, \$14248\, \$12177\, 
               \$10819\, \$13351\, \$13808\, \$15092\, \$10833\, \$12292\, 
               \$11486\, \$14841\, \$15063\, \$14022\, \$10915\, \$12106\, 
               \$13409\, \$10754\, \$15586\, \$14356\, \$13698\, \$15005\, 
               \$12681\, \$11906\, \$15422\, \$12472\, \$15401\, \$11968\, 
               \$10914\, \$11379\, \$14130\, \$12349\, \$14193\, \$11099\, 
               \$11731\, \$10741\, \$14557\, \$12350\, \$11739\, \$12100\, 
               \$10758\, \$12546\, \$12538\, \$11331\, \$12780\, \$14135\, 
               \$14351\, \$11810\, \$12227\, \$13072\, \$14537\, \$15565\, 
               \$13400\, \$13722\, \$12673\, \$14243\, \$12772\, \$10898\, 
               \$12588\, \$13080\, \$12423\, \$12037\ : value(0 to 107) := (others => '0');
      variable \$v6311\, \$12427\, \$14647\, \$11889_i\, \$v5078\, \$v6028\, 
               \$13294\, \$13093\, \$15268\, \$12690\, \$14198\, \$v5714\, 
               \$12289_i\, \$14407\, \$13807\, \$15090_i\, \$v4705\, 
               \$10753\, \$13663_i\, \$14536\, \$v5588\, \$14319_i\, 
               \$12555\, \$15043\, \$v5298\, \$15632\, \$15469\, \$11749\, 
               \$10966_i\, \$11917\, \$15035\, \$v4153\, \$15074\, 
               \$13850_i\, \$15648\, \$v4624\, \$v4708\, \$12884\, 
               \$15128_i\, \$13743_i\, \$v3368\, \$11338\, \$v6141\, 
               \$12829_a\, \$12718_a\, \$v5583\, \$10757\, \$15477\, 
               \$12436\, \$14058_i\, \$v4080\, \$12989\, \$v4962\, \$15644\, 
               \$11222\, \$v5241\, \$10826\, \$v4091\, \$12550\, \$13746\, 
               \$15595_i\, \$15678\, \$11534\, \$13225\, \$10896\, \$v3516\, 
               \$11576\, \$v3655\, \$v6248\, \$v5501\, \$14125_i\, \$v3966\, 
               \$v5898\, \$v5375\, \$10913_i\, \$10792\, \$v5882\, 
               \$14271_i\, \$13783_i\, \$13089\, \$v6647\, \$v3591\, 
               \$14012_i\, \$12039\, \$13399\, \$14655\, \$11420_i\, 
               \$11032_i\, \$v6573\, \$v3981\, \$12604_j\, \$14666\, 
               \$v3683\, \$v6079\, \$v6345\, \$v4883\, \$11218\, \$14192\, 
               \$v6980\, \$v3412\, \$11826\, \$v5591\, \$11504_i\, 
               \$13443_i\, \$13098\, \$15470\, \$12304\, \$v3470\, \$12991\, 
               \$14651\, \$13769_i\, \$13382_i\, \$14728\, \$15594_j\, 
               \$v6577\, \$v4720\, \$11267_i\, \$12291\, \$11466_i\, 
               \$v5561\, \$11668\, \$15628\, \$13684_i\, \$11670\, \$12793\, 
               \$12176\, \$15391_len_aux3143348_result\, \$15131\, \$12308\, 
               \$11594\, \$14642\, \$v6054\, \$v3477\, \$14445_i\, \$11666\, 
               \$v4884\, \$15488\, \$12971\, \$12173\, \$15342\, \$12605_i\, 
               \$11944_i\, \$12384_i\, \$11627_i\, \$10737\, \$13598\, 
               \$15630_i\, \$v5579\, \$v4694\, \$v6140\, \$11293_i\, 
               \$11228_i\, \$v4403\, \$12691_i\, \$v6526\, \$13545_i\, 
               \$15434_j\, \$v4398\, \$12599_i\, \$v5336\, \$15598_j\, 
               \$v3458\, \$v3504\, \$15473\, \$v4423\, \$v3493\, \$v5709\, 
               \$v3807\, \$11708\, \$12616_j\, \$12670_i\, \$13872_j\, 
               \$v4698\, \$v5146\, \$12776\, \$10765\, \$11657\, \$13595_i\, 
               \$11738\, \$11667_i\, \$v4270\, \$15319\, \$v3848\, \$11819\, 
               \$13837\, \$12984\, \$14405_i\, \$13869_i\, \$15262\, 
               \$v3580\, \$12889\, \$15457\, \$11134_i\, \$v6578\, \$v5694\, 
               \$14541\, \$13028_b\, \$10893_i\, \$14472_i\, \$11971\, 
               \$v4217\, \$12122\, \$v4449\, \$11972_i\, \$v5748\, \$v5259\, 
               \$13665\, \$11675\, \$v6330\, \$v6236\, \$14936\, \$12053\, 
               \$15760_i\, \$15306\, \$10767_j\, \$v5832\, \$12607_j\, 
               \$11280_i\, \$12225_i\, \$12190\, \$15298\, \$11213\, 
               \$v6352\, \$11433_i\, \$v3667\, \$v4750\, \$15313\, \$14415\, 
               \$v6901\, \$14837\, \$15611_i\, \$12035\, \$13482_i\, 
               \$14595_i\, \$12110_i\, \$v4684\, \$14211_i\, \$v5337\, 
               \$11905\, \$11596\, \$v6441\, \$v3417\, \$11713\, \$v4589\, 
               \$14681_i\, \$v4973\, \$14658\, \$v5633\, \$v6766\, \$v3717\, 
               \$12879\, \$10766\, \$12261_i\, \$v4679\, \$11406_i\, 
               \$15613_i\, \$15796\, \$13177\, \$10979_i\, \$11665\, 
               \$13626_i\, \$v6897\, \$11787_i\, \$12976\, \$v5289\, 
               \$11655_i\, \$v5799\, \$v3565\, \$13234\, \$14306\, 
               \$13291_i\, \$14079\, \$v5121\, \$12431\, \$14722\, 
               \$15129_i\, \$12083_i\, \$12433_i\, \$15261\, \$14972\, 
               \$14409\, \$v6066\, \$v6584\, \$11147_i\, \$v3465\, \$v4885\, 
               \$12104\, \$15465\, \$v5873\, \$v4438\, \$v6809\, \$13829_i\, 
               \$14580_i\, \$15763_j\, \$v3577\, \$12414\, \$14763_i\, 
               \$v5468\, \$v4609\, \$11730\, \$11321_i\, \$14185_i\, 
               \$13128_b\, \$12614_i\, \$13985_i\, \$12113\, \$12855_i\, 
               \$15431_i\, \$14390_i\, \$v5730\, \$12299\, \$v6605\, 
               \$12309\, \$12993\, \$14158_i\, \$v5349\, \$15506\, \$15324\, 
               \$v3992\, \$14458_i\, \$15471_i\, \$15629\, \$11966\, 
               \$11520_i\, \$14284_i\, \$12313\, \$14705_i\, \$12041_i\, 
               \$v5043\, \$13868_j\, \$12545\, \$v4688\, \$v6261\, \$v6117\, 
               \$12928_b\, \$v5269\, \$14540\, \$12788\, \$15137\, \$v5397\, 
               \$v3894\, \$10842\, \$v5954\, \$11327\, \$14834_i\, 
               \$12556_i\, \$11172_i\, \$15724_len_aux3143361_result\, 
               \$v5810\, \$13741\, \$11236\, \$13129_a\, \$10731\, \$11803\, 
               \$12790_i\, \$12494_i\, \$v5370\, \$15033\, \$v5157\, 
               \$12990_i\, \$v5382\, \$11065_i\, \$11756\, \$14858_i\, 
               \$11006_i\, \$v3592\, \$v6916\, \$15788_get_int268_result\, 
               \$13155_i\, \$14839\, \$15314\, \$v5823\, \$v4805\, \$v6737\, 
               \$11903_i\, \$11571\, \$v4680\, \$v4988\, \$13178_i\, 
               \$v5120\, \$12685\, \$14072_i\, \$13415\, \$12955_i\, 
               \$v4695\, \$v3637\, \$12348_i\, \$13606\, \$10749\, 
               \$12828_b\, \$v5609\, \$12755_i\, \$15293\, \$13972\, 
               \$14650\, \$11121_i\, \$15034_i\, \$15141\, \$15702\, 
               \$v5052\, \$10740\, \$13744\, \$14603\, \$v4596\, 
               \$15555_len_aux3143354_result\, \$15640\, \$13640_i\, 
               \$11748_i\, \$11812\, \$13999_i\, \$12888\, \$14772\, 
               \$v5515\, \$14719_i\, \$15186_i\, \$13718_i\, \$13600_i\, 
               \$12471_i\, \$15673\, \$15032\, \$v3486\, \$v4830\, 
               \$14720_i\, \$11482_i\, \$11560_i\, \$v4804\, \$15454\, 
               \$v4637\, \$12186\, \$14892_i\, \$v4281\, \$12185\, 
               \$12608_i\, \$v3705\, \$14912\, \$12798\, \$v5965\, 
               \$15263_i\, \$11558\, \$v4803\, \$12248_i\, \$12311\, 
               \$v3388\, \$12610_j\, \$v4685\, \$12398_i\, \$v5861\, 
               \$12559\, \$13408\, \$15636\, \$11303\, \$15294\, \$v6380\, 
               \$v6592\, \$12030\, \$14795_i\, \$15479_i\, \$v3374\, 
               \$12876\, \$14404_i\, \$14770\, \$v3674\, \$12042\, 
               \$13529_i\, \$v5970\, \$11848\, \$v5628\, \$v4228\, \$12893\, 
               \$11821\, \$v5772\, \$13252_c\, \$12040\, \$12296\, \$v6483\, 
               \$13404\, \$13495_i\, \$15463_i\, \$13071\, \$15114_i\, 
               \$v6851\, \$v5850\, \$11910\, \$v5122\, \$v5504\, \$12869_i\, 
               \$10827\, \$12629_i\, \$v5587\, \$12979\, \$v4356\, \$15255\, 
               \$v6808\, \$14112_i\, \$v4815\, \$15534\, \$14797\, 
               \$15447_i\, \$13076\, \$10853\, \$12890_i\, \$15637\, 
               \$15305\, \$10734\, \$15478\, \$12097_i\, \$15696\, 
               \$14346_i\, \$15782_i\, \$v4999\, \$v6747\, \$v5612\, 
               \$12188\, \$12275_i\, \$10813\, \$v5990\, \$15481\, \$v6043\, 
               \$11294_i\, \$v4635\, \$15067\, \$15797\, \$11185_i\, 
               \$11808\, \$v5598\, \$13029_a\, \$13742\, \$v4345\, \$v4104\, 
               \$13091\, \$13278_i\, \$15764_i\, \$11801_i\, \$v5635\, 
               \$12891\, \$11539\, \$v4503\, \$11518_i\, \$11221\, 
               \$10940_i\, \$12521_i\, \$11568_i\, \$v6581\, \$11081_i\, 
               \$v4292\, \$v4410\, \$10762\, \$12542\, \$13368_i\, \$13176\, 
               \$v3702\, \$v6755\, \$14665\, \$v5322\, \$11984\, \$13459_i\, 
               \$11084\, \$v4806\, \$v4964\, \$15317\, \$v5277\, \$v6600\, 
               \$12099\, \$14654\, \$13088\, \$12565\, \$15265\, \$14597\, 
               \$v5412\, \$14799\, \$13812\, \$v6059\, \$12181\, \$15307_i\, 
               \$15455\, \$13186\, \$v3694\, \$v4164\, \$v5627\, \$13292_i\, 
               \$11846_i\, \$15483\, \$13229\, \$v4038\, \$12109\, 
               \$12584_j\, \$11818_i\, \$11925\, \$10720\, \$12108\, 
               \$13831\, \$13864_i\, \$15365\, \$11854\, \$v6527\, \$v3391\, 
               \$v6905\, \$11485\, \$14171_i\, \$v3396\, \$v6299\, \$13599\, 
               \$v3909\, \$v5041\, \$v4735\, \$12602_i\, \$12656_i\, 
               \$13169_i\, \$11915\, \$14609\, \$v5584\, \$v5947\, \$v5067\, 
               \$12779\, \$15309\, \$11845\, \$13227\, \$v5131\, \$15075\, 
               \$v5248\, \$12166_i\, \$13347_i\, \$11468_i\, \$14498\, 
               \$v5325\, \$12998\, \$v4496\, \$v4531\, \$15430_j\, 
               \$13886_i\, \$v4102\, \$v3377\, \$12434\, \$15780_i\, 
               \$12028_i\, \$10761\, \$11706_i\, \$10811\, \$11975\, 
               \$v5476\, \$v6889\, \$v5342\, \$11562\, \$12195\, \$v6379\, 
               \$v6565\, \$13613\, \$11330\, \$v4713\, \$15025_i\, 
               \$15638_i\, \$15347\, \$12554\, \$13581_i\, \$11751\, 
               \$15315_i\, \$10763_i\, \$11364_i\, \$15754_i\, \$15511\, 
               \$v5262\, \$v5897\, \$12929_a\, \$15621\, \$13313_i\, 
               \$v6908\, \$14939_get_int268_result\, \$v3424\, \$11550\, 
               \$v6928\, \$v6744\, \$v6902\, \$11816\, \$v5811\, \$13865_i\, 
               \$13084\, \$v4683\, \$13090_i\, \$12371_i\, \$12642_i\, 
               \$11555\, \$12898\, \$v6927\, \$14085\, \$11491\, \$11859\, 
               \$v5042\, \$v5781\, \$14768_i\, \$v6690\, \$13923\, \$v4920\, 
               \$12601_j\, \$v4636\, \$12694\, \$14911\, \$15645\, 
               \$11641_i\, \$v3501\, \$10797_i\, \$11067_i\, \$12310_i\, 
               \$v5816\, \$v3634\, \$11569\, \$13645\, \$v4841\, \$v6225\, 
               \$15299_i\, \$v6898\, \$12717_b\, \$11566\, \$v4704\, 
               \$12613_j\, \$13428_i\, \$13055_i\, \$11547\, \$12537\, 
               \$12412_i\, \$14499\, \$v6741\, \$v4909\, \$13226_i\, 
               \$14897_get_int268_result\, \$11919\, \$11916_i\, \$15622\, 
               \$11351_i\, \$13442_i\, \$13601\, \$13179\, \$11296\, 
               \$12422\, \$v5765\, \$v5199\, \$13603\, \$14640_i\, \$v6595\, 
               \$11559\, \$v6129\, \$v6183\, \$v6740\, \$13069_i\, \$v5977\, 
               \$11844\, \$15301\, \$v5697\, \$15172_i\, \$12969_i\, 
               \$14949_x\, \$13181\, \$v6648\, \$15591_i\, \$14594_i\, 
               \$13756\, \$11970\, \$v3442\, \$13220\, \$10880_i\, 
               \$15646_i\, \$v5488\, \$15529\, \$15585_i\, \$15421_i\, 
               \$v5708\, \$12111\, \$13942\, \$12680\, \$14766_i\, 
               \$11098_i\, \$12583_i\, \$12771\, \$11542\, \$v5796\, 
               \$11743\, \$14225_i\, \$11232\, \$14991_i\, \$v5866\, 
               \$v5415\, \$v6484\, \$12014_i\, \$v5469\, \$v6574\, \$15274\, 
               \$v5426\, \$v6241\, \$15370\, \$13224\, \$12535_i\, 
               \$11019_i\, \$12769_i\, \$15070\, \$v3403\, \$14913_x\, 
               \$11746\, \$12791\, \$v3920\, \$13739_i\, \$v5564\, 
               \$15427_i\, \$13966\, \$v3720\, \$15037\, \$12692\, 
               \$15449_i\, \$v4584\, \$v5270\, \$13445\, \$12611_i\, 
               \$14298_i\, \$11567\, \$15767_j\, \$12441\, \$11662\, 
               \$v4894\, \$v4334\, \$12168\, \$12677\, \$14732\, \$11959_i\, 
               \$14948\, \$13568_i\, \$v4146\, \$11187_i\, \$13749\, 
               \$15650\, \$v4963\, \$12557\, \$14045_i\, \$10867_i\, 
               \$v5944\, \$10736\, \$13816\, \$15256\, \$v4761\, \$v4542\, 
               \$v6736\, \$11961\, \$12784\, \$14777\, \$14377_i\, \$v4491\, 
               \$v3822\, \$v4516\, \$14947\, \$10953_i\, \$14661\, \$10717\, 
               \$v6318\, \$11747\, \$12988\, \$12187_i\, \$12152_i\, 
               \$v6728\, \$12871\, \$11298\, \$14238_i\, \$12689\, \$13079\, 
               \$v5760\, \$11378_i\, \$v5721\, \$v3437\, \$11817\, \$v5847\, 
               \$v5759\, \$13788\, \$15462\, \$14098_i\, \$14803\, \$12044\, 
               \$v5358\, \$13215\, \$11230\, \$14500_x\, \$10838_nargs\, 
               \$13913_i\, \$11735\, \$v3449\, \$v5745\, \$v3369\, 
               \$14333_i\, \$14300\, \$v4103\, \$12672\, \$v3837\, \$12789\, 
               \$15062\, \$11973\, \$v3662\, \$v4206\, \$12318\, \$10810\, 
               \$v3523\, \$12507_i\, \$15655\, \$12432\, \$v5634\, \$11914\, 
               \$12419\, \$12699\, \$v3652\, \$15296\, \$14556_i\, 
               \$15798_x\, \$11728_i\ : value(0 to 31) := (others => '0');
      variable \$$10695_limit_ptr_take\ : value(0 to 0) := "0";
      variable \$$10696_ram_ptr_take\ : value(0 to 0) := "0";
      variable \$$10697_stack_ptr_take\ : value(0 to 0) := "0";
      variable \$$10698_heap_ptr_take\ : value(0 to 0) := "0";
      variable \$$10699_symtbl_ptr_take\ : value(0 to 0) := "0";
      variable \$$10700_pc_ptr_take\ : value(0 to 0) := "0";
      variable \$$10701_pos_ptr_take\ : value(0 to 0) := "0";
      variable \$$10702_brk_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$15391_len_aux3143348_arg\); default_zero(\$v6130\); 
          default_zero(\$v6642\); default_zero(\$v4211\); 
          default_zero(\$11728_i\); default_zero(\$15798_x\); 
          default_zero(\$14556_i\); default_zero(\$v6071\); 
          default_zero(\$12037\); default_zero(\$v3571\); 
          default_zero(\$v5232\); default_zero(\$12423\); 
          default_zero(\$15296\); default_zero(\$v3718\); 
          default_zero(\$v3652\); default_zero(\$12699\); 
          default_zero(\$v4604\); default_zero(\$12419\); 
          default_zero(\$11914\); default_zero(\$v5634\); 
          default_zero(\$v5442\); default_zero(\$12432\); 
          default_zero(\$v4325\); default_zero(\$15655\); 
          default_zero(\$v6512\); default_zero(\$12507_i\); 
          default_zero(\$v3523\); default_zero(\$v6070\); 
          default_zero(\$10810\); default_zero(\$v4079\); 
          default_zero(\$v4874\); default_zero(\$v4120\); 
          default_zero(\$v5152\); default_zero(\$12318\); 
          default_zero(\$13689_list_tail2653276_arg\); 
          default_zero(\$v4206\); default_zero(\$v4703\); 
          default_zero(\$v3662\); default_zero(\$v4814\); 
          default_zero(\$v4710\); default_zero(\$11973\); 
          default_zero(\$v5458\); default_zero(\$15062\); 
          default_zero(\$v4781\); default_zero(\$12789\); 
          default_zero(\$v4610\); default_zero(\$v3837\); 
          default_zero(\$12672\); default_zero(\$v5282\); 
          default_zero(\$v4103\); default_zero(\$v3824\); 
          default_zero(\$14300\); default_zero(\$14333_i\); 
          default_zero(\$v3369\); default_zero(\$v3402\); 
          default_zero(\$v6240\); default_zero(\$11564_r\); 
          default_zero(\$v5616\); default_zero(\$v4904\); 
          default_zero(\$v5745\); default_zero(\$v3449\); 
          default_zero(\$v6128\); default_zero(\$v6199\); 
          default_zero(\$11735\); default_zero(\$v5592\); 
          default_zero(\$v4760\); default_zero(\$13913_i\); 
          default_zero(\$10838_nargs\); default_zero(\$14500_x\); 
          default_zero(\$v4749\); default_zero(\$v4486\); 
          default_zero(\$v3462\); default_zero(\$v5369\); 
          default_zero(\$v4741\); default_zero(\$14659\); 
          default_zero(\$11230\); default_zero(\$13215\); 
          default_zero(\$v5358\); default_zero(\$v5414\); 
          default_zero(\$v5945\); default_zero(\$12044\); 
          default_zero(\$14803\); default_zero(\$v4725\); 
          default_zero(\$14098_i\); default_zero(\$15462\); 
          default_zero(\$v4437\); default_zero(\$v4050\); 
          default_zero(\$v5752\); default_zero(\$v4084\); 
          default_zero(\$13788\); default_zero(\$v5407\); 
          default_zero(\$v5759\); default_zero(\$v6855\); 
          default_zero(\$v5836\); default_zero(\$v5847\); 
          default_zero(\$11817\); default_zero(\$v3437\); 
          default_zero(\$v5703\); default_zero(\$v3382\); 
          default_zero(\$v5721\); default_zero(\$11378_i\); 
          default_zero(\$v5952\); default_zero(\$v5935\); 
          default_zero(\$v5760\); default_zero(\$v5137\); 
          default_zero(\$v5931\); default_zero(\$v3453\); 
          default_zero(\$v3798\); default_zero(\$13079\); 
          default_zero(\$v3919\); default_zero(\$12689\); 
          default_zero(\$v5019\); default_zero(\$v6967\); 
          default_zero(\$v4300\); default_zero(\$14238_i\); 
          default_zero(\$v4416\); default_zero(\$11298\); 
          default_zero(\$v6027\); default_zero(\$v6078\); 
          default_zero(\$12871\); default_zero(\$v6728\); 
          default_zero(\$v6500\); default_zero(\$v4603\); 
          default_zero(\$v6496\); default_zero(\$v6894\); 
          default_zero(\$v6470\); default_zero(\$v5610\); 
          default_zero(\$v4952\); default_zero(\$13446\); 
          default_zero(\$12152_i\); default_zero(\$12187_i\); 
          default_zero(\$12988\); default_zero(\$v4029\); 
          default_zero(\$v4692\); default_zero(\$13080\); 
          default_zero(\$12588\); default_zero(\$11747\); 
          default_zero(\$v6599\); default_zero(\$v6318\); 
          default_zero(\$v5364\); default_zero(\$10717\); 
          default_zero(\$14661\); default_zero(\$10953_i\); 
          default_zero(\$14947\); default_zero(\$v5777\); 
          default_zero(\$v4516\); default_zero(\$v3822\); 
          default_zero(\$v3508\); default_zero(\$v4004\); 
          default_zero(\$v4491\); default_zero(\$v4054\); 
          default_zero(\$14377_i\); default_zero(\$14777\); 
          default_zero(\$12784\); default_zero(\$v4734\); 
          default_zero(\$10898\); default_zero(\$v5655\); 
          default_zero(\$v5838\); default_zero(\$11961\); 
          default_zero(\$v3699\); default_zero(\$v4351\); 
          default_zero(\$v6736\); default_zero(\$v5604\); 
          default_zero(\$12772\); default_zero(\$v4542\); 
          default_zero(\$v6508\); default_zero(\$v4761\); 
          default_zero(\$v6591\); default_zero(\$15256\); 
          default_zero(\$v6095\); default_zero(\$13816\); 
          default_zero(\$v4276\); default_zero(\$10736\); 
          default_zero(\$v5582\); default_zero(\$v6211\); 
          default_zero(\$v3967\); default_zero(\$v4136\); 
          default_zero(\$v5944\); default_zero(\$v4116\); 
          default_zero(\$10867_i\); default_zero(\$14243\); 
          default_zero(\$v4280\); default_zero(\$v4417\); 
          default_zero(\$14045_i\); default_zero(\$v6732\); 
          default_zero(\$12557\); default_zero(\$v4963\); 
          default_zero(\$v3847\); default_zero(\$v3957\); 
          default_zero(\$v5639\); default_zero(\$15650\); 
          default_zero(\$13749\); default_zero(\$11187_i\); 
          default_zero(\$v3876\); default_zero(\$v4146\); 
          default_zero(\$13568_i\); default_zero(\$v6058\); 
          default_zero(\$v4674\); default_zero(\$v5250\); 
          default_zero(\$14948\); default_zero(\$v6323\); 
          default_zero(\$11959_i\); default_zero(\$14732\); 
          default_zero(\$12677\); default_zero(\$12168\); 
          default_zero(\$v3604\); default_zero(\$v4334\); 
          default_zero(\$v5958\); default_zero(\$v4894\); 
          default_zero(\$12673\); default_zero(\$11662\); 
          default_zero(\$12441\); default_zero(\$15767_j\); 
          default_zero(\$11567\); default_zero(\$v5430\); 
          default_zero(\$v3629\); default_zero(\$v6513\); 
          default_zero(\$13722\); default_zero(\$14298_i\); 
          default_zero(\$12611_i\); default_zero(\$v3809\); 
          default_zero(\$v5514\); default_zero(\$v4148\); 
          default_zero(\$v4634\); default_zero(\$13445\); 
          default_zero(\$v6723\); default_zero(\$v4097\); 
          default_zero(\$v6746\); default_zero(\$v5270\); 
          default_zero(\$v4584\); 
          default_zero(\$13500_list_tail2653266_arg\); 
          default_zero(\$v6038\); default_zero(\$v4711\); 
          default_zero(\$v5735\); default_zero(\$15449_i\); 
          default_zero(\$12692\); default_zero(\$v6733\); 
          default_zero(\$14667_new_rib\); default_zero(\$15037\); 
          default_zero(\$v4641\); default_zero(\$v3720\); 
          default_zero(\$v4393\); default_zero(\$13966\); 
          default_zero(\$v4433\); default_zero(\$v6551\); 
          default_zero(\$13400\); default_zero(\$15565\); 
          default_zero(\$v3698\); default_zero(\$v4928\); 
          default_zero(\$15427_i\); default_zero(\$15311_end_rib\); 
          default_zero(\$v5284\); default_zero(\$v5564\); 
          default_zero(\$13739_i\); default_zero(\$v3920\); 
          default_zero(\$12791\); default_zero(\$11746\); 
          default_zero(\$v5519\); default_zero(\$v5046\); 
          default_zero(\$14913_x\); default_zero(\$v3403\); 
          default_zero(\$v6131\); default_zero(\$15070\); 
          default_zero(\$v3904\); default_zero(\$v6914\); 
          default_zero(\$v5247\); default_zero(\$v5420\); 
          default_zero(\$12769_i\); default_zero(\$14537\); 
          default_zero(\$11019_i\); default_zero(\$v5027\); 
          default_zero(\$v5069\); default_zero(\$10840\); 
          default_zero(\$v5860\); default_zero(\$12036\); 
          default_zero(\$v4414\); default_zero(\$v3641\); 
          default_zero(\$v3390\); default_zero(\$12535_i\); 
          default_zero(\$13224\); default_zero(\$15370\); 
          default_zero(\$v6241\); default_zero(\$v5426\); 
          default_zero(\$v5539\); default_zero(\$v6593\); 
          default_zero(\$v6884\); default_zero(\$v4425\); 
          default_zero(\$15274\); default_zero(\$v5870\); 
          default_zero(\$v6461\); default_zero(\$v6574\); 
          default_zero(\$v5469\); default_zero(\$15267\); 
          default_zero(\$v4574\); default_zero(\$v4661\); 
          default_zero(\$v5203\); default_zero(\$12014_i\); 
          default_zero(\$v4409\); default_zero(\$v3635\); 
          default_zero(\$v6484\); default_zero(\$v5415\); 
          default_zero(\$v4699\); default_zero(\$v6428\); 
          default_zero(\$v5123\); default_zero(\$v5866\); 
          default_zero(\$v5951\); default_zero(\$14991_i\); 
          default_zero(\$12885_y\); default_zero(\$11232\); 
          default_zero(\$15724_len_aux3143361_arg\); default_zero(\$v5148\); 
          default_zero(\$v5815\); default_zero(\$14225_i\); 
          default_zero(\$11743\); default_zero(\$v4798\); 
          default_zero(\$v5846\); default_zero(\$v3987\); 
          default_zero(\$v6986\); default_zero(\$v6702\); 
          default_zero(\$v4248\); default_zero(\$v5796\); 
          default_zero(\$v6277\); default_zero(\$11542\); 
          default_zero(\$12771\); default_zero(\$v5985\); 
          default_zero(\$v4756\); default_zero(\$12583_i\); 
          default_zero(\$v5795\); default_zero(\$v4453\); 
          default_zero(\$11098_i\); default_zero(\$14766_i\); 
          default_zero(\$11196_loop2913158_result\); default_zero(\$v5132\); 
          default_zero(\$v6913\); default_zero(\$12680\); 
          default_zero(\$13942\); default_zero(\$v4541\); 
          default_zero(\$v6344\); default_zero(\$v4975\); 
          default_zero(\$12111\); default_zero(\$v6896\); 
          default_zero(\$v6906\); default_zero(\$v5647\); 
          default_zero(\$v5357\); default_zero(\$v5708\); 
          default_zero(\$15421_i\); default_zero(\$15585_i\); 
          default_zero(\$15529\); default_zero(\$v5488\); 
          default_zero(\$v4368\); default_zero(\$v4184\); 
          default_zero(\$v4895\); default_zero(\$v5580\); 
          default_zero(\$v4067\); default_zero(\$15646_i\); 
          default_zero(\$v4893\); default_zero(\$v4924\); 
          default_zero(\$10880_i\); default_zero(\$v5031\); 
          default_zero(\$v4188\); default_zero(\$v5161\); 
          default_zero(\$13220\); default_zero(\$v5450\); 
          default_zero(\$v4112\); default_zero(\$v3996\); 
          default_zero(\$v6753\); default_zero(\$v3442\); 
          default_zero(\$v6482\); default_zero(\$11970\); 
          default_zero(\$13756\); default_zero(\$v5611\); 
          default_zero(\$13072\); default_zero(\$14594_i\); 
          default_zero(\$15591_i\); default_zero(\$v6648\); 
          default_zero(\$v6751\); default_zero(\$v5651\); 
          default_zero(\$13181\); default_zero(\$v5589\); 
          default_zero(\$v4384\); default_zero(\$v6453\); 
          default_zero(\$v6103\); default_zero(\$v3839\); 
          default_zero(\$14949_x\); default_zero(\$v3407\); 
          default_zero(\$12969_i\); default_zero(\$15172_i\); 
          default_zero(\$v6738\); default_zero(\$12227\); 
          default_zero(\$v5697\); default_zero(\$15301\); 
          default_zero(\$11844\); default_zero(\$10818_proc\); 
          default_zero(\$v6034\); default_zero(\$v6065\); 
          default_zero(\$v5977\); default_zero(\$13069_i\); 
          default_zero(\$v4965\); default_zero(\$v5878\); 
          default_zero(\$v3673\); default_zero(\$v6740\); 
          default_zero(\$v6183\); default_zero(\$v6129\); 
          default_zero(\$v5379\); default_zero(\$11810\); 
          default_zero(\$11559\); default_zero(\$v6350\); 
          default_zero(\$v6595\); default_zero(\$14640_i\); 
          default_zero(\$v4500\); default_zero(\$13603\); 
          default_zero(\$14351\); default_zero(\$v6629\); 
          default_zero(\$v4490\); default_zero(\$v4159\); 
          default_zero(\$v5199\); default_zero(\$v4163\); 
          default_zero(\$v5765\); default_zero(\$v5044\); 
          default_zero(\$v3492\); default_zero(\$12422\); 
          default_zero(\$11296\); default_zero(\$v3961\); 
          default_zero(\$v3408\); default_zero(\$v4696\); 
          default_zero(\$13179\); default_zero(\$13601\); 
          default_zero(\$v4619\); default_zero(\$v6761\); 
          default_zero(\$13442_i\); default_zero(\$v4537\); 
          default_zero(\$11351_i\); default_zero(\$15622\); 
          default_zero(\$11916_i\); default_zero(\$11919\); 
          default_zero(\$14897_get_int268_result\); default_zero(\$v4518\); 
          default_zero(\$13226_i\); default_zero(\$v4909\); 
          default_zero(\$v3777\); default_zero(\$v6741\); 
          default_zero(\$v5656\); default_zero(\$14499\); 
          default_zero(\$12412_i\); default_zero(\$14135\); 
          default_zero(\$v4408\); default_zero(\$11323\); 
          default_zero(\$v6656\); default_zero(\$12537\); 
          default_zero(result3362); default_zero(\$v6014\); 
          default_zero(\$v4407\); default_zero(\$v5003\); 
          default_zero(\$11547\); default_zero(\$v3474\); 
          default_zero(\$13055_i\); default_zero(\$v5398\); 
          default_zero(\$13428_i\); default_zero(\$12613_j\); 
          default_zero(\$v4176\); default_zero(\$v6044\); 
          default_zero(\$v4704\); default_zero(\$11566\); 
          default_zero(\$12717_b\); default_zero(\$v3579\); 
          default_zero(\$v6898\); default_zero(\$15299_i\); 
          default_zero(\$v3666\); default_zero(\$v6225\); 
          default_zero(\$v4841\); default_zero(\$v6121\); 
          default_zero(\$13645\); default_zero(\$v3625\); 
          default_zero(\$v3794\); default_zero(\$v5467\); 
          default_zero(\$v4886\); default_zero(\$v3410\); 
          default_zero(\$v6594\); default_zero(\$v6207\); 
          default_zero(\$v6971\); default_zero(\$v5769\); 
          default_zero(\$11569\); default_zero(\$11540_x\); 
          default_zero(\$v3634\); default_zero(\$v3968\); 
          default_zero(\$v5419\); default_zero(\$12886\); 
          default_zero(\$v5816\); default_zero(\$12780\); 
          default_zero(\$12310_i\); default_zero(\$v4201\); 
          default_zero(\$11067_i\); default_zero(\$10797_i\); 
          default_zero(\$v4389\); default_zero(\$v4807\); 
          default_zero(\$v6265\); default_zero(\$v5608\); 
          default_zero(\$v3501\); default_zero(\$v4071\); 
          default_zero(\$11331\); default_zero(\$v4682\); 
          default_zero(\$v4338\); default_zero(\$v5599\); 
          default_zero(\$11641_i\); default_zero(\$v3802\); 
          default_zero(\$v4998\); default_zero(\$15645\); 
          default_zero(\$14911\); default_zero(\$v3785\); 
          default_zero(\$v5994\); default_zero(\$v6049\); 
          default_zero(\$v5281\); default_zero(\$v4282\); 
          default_zero(\$12694\); default_zero(\$v4636\); 
          default_zero(\$v5574\); default_zero(\$v5015\); 
          default_zero(\$v4062\); default_zero(\$v4429\); 
          default_zero(\$12601_j\); default_zero(\$v4418\); 
          default_zero(\$v6042\); default_zero(\$14973\); 
          default_zero(\$v5082\); default_zero(\$v4920\); 
          default_zero(\$13923\); default_zero(\$v5227\); 
          default_zero(\$v3761\); default_zero(\$v3642\); 
          default_zero(\$v6690\); default_zero(\$v6765\); 
          default_zero(\$14768_i\); default_zero(\$v5781\); 
          default_zero(\$v6900\); default_zero(\$v5042\); 
          default_zero(\$12538\); default_zero(\$v6543\); 
          default_zero(\$v5086\); default_zero(\$13174\); 
          default_zero(\$11859\); default_zero(\$11491\); 
          default_zero(\$v4593\); default_zero(\$14085\); 
          default_zero(\$12546\); default_zero(\$v4865\); 
          default_zero(\$v6927\); default_zero(\$10758\); 
          default_zero(\$12898\); default_zero(\$12100\); 
          default_zero(\$11555\); default_zero(\$v3821\); 
          default_zero(\$v6743\); default_zero(\$12642_i\); 
          default_zero(\$v5054\); default_zero(\$v6742\); 
          default_zero(\$11739\); default_zero(\$v4324\); 
          default_zero(\$v4440\); default_zero(\$v3823\); 
          default_zero(\$12371_i\); default_zero(\$13090_i\); 
          default_zero(\$v7020\); default_zero(\$v6786\); 
          default_zero(\$v4683\); default_zero(\$13084\); 
          default_zero(\$13865_i\); default_zero(\$v4196\); 
          default_zero(\$v5487\); default_zero(\$v5811\); 
          default_zero(\$12350\); default_zero(\$v3651\); 
          default_zero(\$v4376\); default_zero(\$v6547\); 
          default_zero(\$11816\); default_zero(\$v6902\); 
          default_zero(\$v5446\); default_zero(\$v6087\); 
          default_zero(\$v6744\); default_zero(\$v6928\); 
          default_zero(\$11550\); default_zero(\$v3424\); 
          default_zero(\$v5295\); default_zero(\$v4882\); 
          default_zero(\$14939_get_int268_result\); default_zero(\$v6908\); 
          default_zero(\$13313_i\); default_zero(\$v4615\); 
          default_zero(\$15621\); default_zero(\$v6023\); 
          default_zero(\$v5309\); default_zero(\$v3509\); 
          default_zero(\$12929_a\); default_zero(\$v5897\); 
          default_zero(\$v5262\); default_zero(\$15634_str_rib\); 
          default_zero(\$15511\); default_zero(\$15754_i\); 
          default_zero(\$v4887\); default_zero(\$11364_i\); 
          default_zero(\$10763_i\); default_zero(\$v4594\); 
          default_zero(\$15315_i\); default_zero(\$v3654\); 
          default_zero(\$v6790\); default_zero(\$v5066\); 
          default_zero(\$v6329\); default_zero(\$v5425\); 
          default_zero(\$v4700\); default_zero(\$11036_loop3073149_arg\); 
          default_zero(\$v4940\); default_zero(\$v6899\); 
          default_zero(\$v6694\); default_zero(\$11751\); 
          default_zero(\$v6356\); default_zero(\$13581_i\); 
          default_zero(\$12554\); default_zero(\$15347\); 
          default_zero(\$15638_i\); default_zero(\$15025_i\); 
          default_zero(\$v4713\); default_zero(\$v3389\); 
          default_zero(\$v4821\); default_zero(\$v5249\); 
          default_zero(\$11330\); default_zero(\$v5664\); 
          default_zero(\$13613\); default_zero(\$v6734\); 
          default_zero(\$v6565\); default_zero(\$v6880\); 
          default_zero(\$v6829\); default_zero(\$v6379\); 
          default_zero(\$v3518\); default_zero(\$12195\); 
          default_zero(\$14557\); default_zero(\$12174_x\); 
          default_zero(\$10741\); default_zero(\$v3781\); 
          default_zero(\$v3464\); default_zero(\$v5964\); 
          default_zero(\$11562\); default_zero(\$v3517\); 
          default_zero(\$v5386\); default_zero(\$v5342\); 
          default_zero(\$v6889\); default_zero(\$v5476\); 
          default_zero(\$11975\); default_zero(\$10811\); 
          default_zero(\$v4793\); default_zero(\$v5622\); 
          default_zero(\$v4972\); default_zero(\$11731\); 
          default_zero(\$11706_i\); default_zero(\$v5254\); 
          default_zero(\$v3482\); default_zero(\$10761\); 
          default_zero(\$v6588\); default_zero(\$v6256\); 
          default_zero(\$11099\); default_zero(\$v5707\); 
          default_zero(\$v4736\); default_zero(\$12028_i\); 
          default_zero(\$14193\); default_zero(\$v6589\); 
          default_zero(\$v6053\); default_zero(\$v3421\); 
          default_zero(\$v3590\); default_zero(\$v6719\); 
          default_zero(\$14996_list_tail2653334_result\); 
          default_zero(\$v5998\); default_zero(\$v4832\); 
          default_zero(\$15780_i\); default_zero(\$v4562\); 
          default_zero(\$v5855\); default_zero(\$12434\); 
          default_zero(\$v4132\); default_zero(\$v5145\); 
          default_zero(\$v3377\); default_zero(\$v5304\); 
          default_zero(\$v4773\); default_zero(\$v6917\); 
          default_zero(\$v4102\); default_zero(\$v6981\); 
          default_zero(\$v5693\); default_zero(\$13886_i\); 
          default_zero(\$v6617\); default_zero(\$15430_j\); 
          default_zero(\$v4274\); default_zero(\$v3564\); 
          default_zero(\$v4948\); default_zero(\$v4531\); 
          default_zero(\$v4496\); default_zero(\$v6247\); 
          default_zero(\$v6474\); default_zero(\$12998\); 
          default_zero(\$v5325\); default_zero(\$v3711\); 
          default_zero(\$v5753\); default_zero(\$14498\); 
          default_zero(\$11468_i\); default_zero(\$13347_i\); 
          default_zero(\$v5865\); default_zero(\$v3881\); 
          default_zero(\$v3576\); default_zero(\$12166_i\); 
          default_zero(\$10778_run286_result\); default_zero(\$v5248\); 
          default_zero(\$15075\); default_zero(\$v6956\); 
          default_zero(\$v6752\); default_zero(\$v5131\); 
          default_zero(\$13227\); default_zero(\$v4873\); 
          default_zero(\$v4689\); default_zero(\$11845\); 
          default_zero(\$v3515\); default_zero(\$v3612\); 
          default_zero(\$v5744\); default_zero(\$v6378\); 
          default_zero(\$v3616\); default_zero(\$15309\); 
          default_zero(\$v5194\); default_zero(\$15642_end_rib\); 
          default_zero(\$v5411\); default_zero(\$v5347\); 
          default_zero(\$12779\); default_zero(\$v5067\); 
          default_zero(\$v4482\); default_zero(\$v4510\); 
          default_zero(\$v5947\); default_zero(\$v5434\); 
          default_zero(\$v4507\); default_zero(\$v4192\); 
          default_zero(\$13814\); default_zero(\$v5584\); 
          default_zero(\$v5023\); default_zero(\$v4501\); 
          default_zero(\$14609\); default_zero(\$v5313\); 
          default_zero(\$v3671\); default_zero(\$v6436\); 
          default_zero(\$v5293\); default_zero(\$v6227\); 
          default_zero(\$11915\); default_zero(\$v3710\); 
          default_zero(\$13169_i\); default_zero(\$12656_i\); 
          default_zero(\$11967\); default_zero(\$14511_loop311_arg\); 
          default_zero(\$11036_loop3073149_result\); default_zero(\$v5185\); 
          default_zero(\$v3556\); default_zero(\$v6531\); 
          default_zero(\$12349\); default_zero(\$12551_y\); 
          default_zero(\$12602_i\); default_zero(\$v4735\); 
          default_zero(\$v5041\); default_zero(\$v3481\); 
          default_zero(\$v4690\); default_zero(\$v3909\); 
          default_zero(\$v6253\); default_zero(\$v6504\); 
          default_zero(\$13599\); default_zero(\$v6907\); 
          default_zero(\$v5296\); default_zero(\$v6299\); 
          default_zero(\$v5689\); default_zero(\$v3396\); 
          default_zero(\$14171_i\); default_zero(\$v6149\); 
          default_zero(\$11485\); default_zero(\$v4719\); 
          default_zero(\$v6677\); default_zero(\$v4240\); 
          default_zero(\$v6905\); default_zero(\$v3391\); 
          default_zero(\$14130\); default_zero(\$v6527\); 
          default_zero(\$v4227\); default_zero(\$v4320\); 
          default_zero(\$v3584\); default_zero(\$v5494\); 
          default_zero(\$11379\); default_zero(\$11854\); 
          default_zero(\$v3982\); default_zero(\$v5389\); 
          default_zero(\$15365\); default_zero(\$v4075\); 
          default_zero(\$v4809\); default_zero(\$v6813\); 
          default_zero(\$13864_i\); default_zero(\$v5094\); 
          default_zero(\$v4312\); default_zero(\$13831\); 
          default_zero(\$v6322\); default_zero(\$v6982\); 
          default_zero(\$v6002\); default_zero(\$12108\); 
          default_zero(\$10720\); default_zero(\$v5543\); 
          default_zero(\$11925\); default_zero(\$11818_i\); 
          default_zero(\$v4461\); default_zero(\$10914\); 
          default_zero(\$12584_j\); default_zero(\$12109\); 
          default_zero(\$v5785\); default_zero(\$v4038\); 
          default_zero(\$11968\); default_zero(\$v6948\); 
          default_zero(\$v5243\); default_zero(\$13229\); 
          default_zero(\$v4066\); default_zero(\$v5849\); 
          default_zero(\$15483\); default_zero(\$11846_i\); 
          default_zero(\$12986\); default_zero(\$v6340\); 
          default_zero(\$v3522\); default_zero(\$13292_i\); 
          default_zero(\$v3423\); default_zero(\$v5627\); 
          default_zero(\$v4164\); default_zero(\$15401\); 
          default_zero(\$v3694\); default_zero(\$v3679\); 
          default_zero(\$13186\); default_zero(\$v5303\); 
          default_zero(\$v3693\); default_zero(\$v3441\); 
          default_zero(\$v6324\); default_zero(\$v4533\); 
          default_zero(\$v3575\); default_zero(\$v5685\); 
          default_zero(\$v6583\); default_zero(\$v5585\); 
          default_zero(\$15455\); default_zero(\$v5960\); 
          default_zero(\$v5459\); default_zero(\$v5181\); 
          default_zero(\$15307_i\); default_zero(\$12181\); 
          default_zero(\$12472\); default_zero(\$v3485\); 
          default_zero(\$10738_main_rib\); default_zero(\$15422\); 
          default_zero(\$v6059\); default_zero(\$v6358\); 
          default_zero(\$v3566\); default_zero(\$v5695\); 
          default_zero(\$13812\); default_zero(\$v5770\); 
          default_zero(\$v5888\); default_zero(\$v6294\); 
          default_zero(\$14799\); default_zero(\$v5412\); 
          default_zero(\$14597\); default_zero(\$v6778\); 
          default_zero(\$v5032\); 
          default_zero(\$13689_list_tail2653276_result\); 
          default_zero(\$v4530\); default_zero(\$15265\); 
          default_zero(\$12565\); default_zero(\$13088\); 
          default_zero(\$v5283\); default_zero(\$v5617\); 
          default_zero(\$14654\); default_zero(\$v4448\); 
          default_zero(\$v4910\); default_zero(\$12099\); 
          default_zero(\$11906\); default_zero(\$v3757\); 
          default_zero(\$v4333\); default_zero(\$v6600\); 
          default_zero(\$v6582\); default_zero(\$v3446\); 
          default_zero(\$v6174\); default_zero(\$v4232\); 
          default_zero(\$v6423\); default_zero(\$v4816\); 
          default_zero(\$v5626\); default_zero(\$v5277\); 
          default_zero(\$15317\); default_zero(\$v4964\); 
          default_zero(\$v4806\); default_zero(\$v3688\); 
          default_zero(\$v6774\); default_zero(\$v3908\); 
          default_zero(\$11084\); default_zero(\$13459_i\); 
          default_zero(\$v5578\); default_zero(\$11984\); 
          default_zero(\$v5362\); default_zero(\$v5322\); 
          default_zero(\$14665\); default_zero(\$v6083\); 
          default_zero(\$v5211\); default_zero(\$v6755\); 
          default_zero(\$v3702\); default_zero(\$v3401\); 
          default_zero(\$13813\); default_zero(\$13176\); 
          default_zero(\$13368_i\); default_zero(\$15399\); 
          default_zero(\$v4730\); default_zero(\$12542\); 
          default_zero(\$v5736\); default_zero(\$v6926\); 
          default_zero(\$10762\); default_zero(\$v4410\); 
          default_zero(\$v6417\); default_zero(\$v3944\); 
          default_zero(\$v6517\); default_zero(\$v3436\); 
          default_zero(\$v3789\); default_zero(\$v6178\); 
          default_zero(\$v4752\); default_zero(\$v4219\); 
          default_zero(\$v4974\); default_zero(\$v3498\); 
          default_zero(\$v5177\); default_zero(\$v4707\); 
          default_zero(\$v4292\); default_zero(\$v6440\); 
          default_zero(\$v3700\); default_zero(\$v3832\); 
          default_zero(\$11081_i\); default_zero(\$v5918\); 
          default_zero(\$v6581\); default_zero(\$11568_i\); 
          default_zero(\$v3948\); default_zero(\$v6895\); 
          default_zero(\$14652_code_proc_rib\); default_zero(\$12521_i\); 
          default_zero(\$v5374\); default_zero(\$12681\); 
          default_zero(\$v3454\); default_zero(\$v5593\); 
          default_zero(\$10940_i\); default_zero(\$v6363\); 
          default_zero(\$v4849\); default_zero(\$11221\); 
          default_zero(\$v6220\); default_zero(\$11518_i\); 
          default_zero(\$v4503\); default_zero(\$v5493\); 
          default_zero(\$v4124\); default_zero(\$15005\); 
          default_zero(\$v5302\); default_zero(\$11539\); 
          default_zero(\$12891\); default_zero(\$v5927\); 
          default_zero(\$13698\); default_zero(\$v6316\); 
          default_zero(\$v3856\); default_zero(\$15732\); 
          default_zero(\$v5635\); default_zero(\$v3608\); 
          default_zero(\$11801_i\); default_zero(\$v3586\); 
          default_zero(\$v3911\); default_zero(\$14356\); 
          default_zero(\$15764_i\); default_zero(\$13278_i\); 
          default_zero(\$13091\); default_zero(\$v4104\); 
          default_zero(\$v4785\); default_zero(\$v4345\); 
          default_zero(\$13742\); default_zero(\$13029_a\); 
          default_zero(\$v5598\); default_zero(\$v3704\); 
          default_zero(\$v4344\); default_zero(\$11808\); 
          default_zero(\$11185_i\); default_zero(\$v6260\); 
          default_zero(\$v4697\); default_zero(\$v4304\); 
          default_zero(\$v4765\); default_zero(\$15797\); 
          default_zero(\$v4649\); default_zero(\$v4316\); 
          default_zero(\$v6698\); default_zero(\$v4223\); 
          default_zero(\$15067\); default_zero(\$v4635\); 
          default_zero(\$11294_i\); default_zero(\$v6043\); 
          default_zero(\$v4968\); default_zero(\$v5820\); 
          default_zero(\$v4686\); default_zero(\$v3885\); 
          default_zero(\$v6842\); default_zero(\$15481\); 
          default_zero(\$v5990\); default_zero(\$v3976\); 
          default_zero(\$10813\); default_zero(\$12275_i\); 
          default_zero(\$15586\); default_zero(\$v6556\); 
          default_zero(\$v5969\); default_zero(\$10754\); 
          default_zero(\$v6195\); default_zero(\$12687\); 
          default_zero(\$12188\); default_zero(\$v3560\); 
          default_zero(\$v5612\); default_zero(\$v6747\); 
          default_zero(\$v5719\); default_zero(\$v4999\); 
          default_zero(\$13409\); default_zero(\$v6331\); 
          default_zero(\$v6169\); default_zero(\$v3680\); 
          default_zero(\$15782_i\); default_zero(\$v6281\); 
          default_zero(\$14346_i\); default_zero(\$v6539\); 
          default_zero(\$15696\); default_zero(\$12097_i\); 
          default_zero(\$v6850\); default_zero(\$15478\); 
          default_zero(\$v3620\); default_zero(\$v6727\); 
          default_zero(\$10734\); default_zero(\$15305\); 
          default_zero(\$15637\); default_zero(\$12890_i\); 
          default_zero(\$v6770\); default_zero(\$12106\); 
          default_zero(\$13221\); default_zero(\$10853\); 
          default_zero(\$13076\); default_zero(\$v4517\); 
          default_zero(\$v5740\); default_zero(\$v3765\); 
          default_zero(\$15447_i\); default_zero(\$14797\); 
          default_zero(\$15534\); default_zero(\$v7006\); 
          default_zero(\$v5879\); default_zero(\$14656_proc_rib\); 
          default_zero(\$v4815\); default_zero(\$v5355\); 
          default_zero(\$14112_i\); default_zero(\$v6808\); 
          default_zero(\$10915\); default_zero(\$v6006\); 
          default_zero(\$v5974\); default_zero(\$v4145\); 
          default_zero(\$v6837\); default_zero(\$12977_x\); 
          default_zero(\$14022\); default_zero(\$v5600\); 
          default_zero(\$15255\); default_zero(\$v5926\); 
          default_zero(\$v4356\); default_zero(\$v3728\); 
          default_zero(\$v4093\); default_zero(\$12979\); 
          default_zero(\$v3880\); default_zero(\$v5587\); 
          default_zero(\$15400\); default_zero(\$12629_i\); 
          default_zero(\$v5804\); default_zero(\$10827\); 
          default_zero(\$v6871\); default_zero(\$12869_i\); 
          default_zero(\$v5842\); default_zero(\$v5267\); 
          default_zero(\$v5527\); default_zero(\$v6757\); 
          default_zero(\$v5258\); default_zero(\$15063\); 
          default_zero(\$v5504\); default_zero(\$v5122\); 
          default_zero(\$v4522\); default_zero(\$11910\); 
          default_zero(\$13318_list_tail2653256_result\); 
          default_zero(\$v5850\); 
          default_zero(\$14996_list_tail2653334_arg\); 
          default_zero(\$13077_x\); default_zero(\$v6851\); 
          default_zero(\$v6018\); default_zero(\$v6888\); 
          default_zero(\$15114_i\); default_zero(\$13071\); 
          default_zero(\$12182_y\); default_zero(\$15463_i\); 
          default_zero(\$v4275\); default_zero(\$13495_i\); 
          default_zero(\$13404\); default_zero(\$14841\); 
          default_zero(\$v5786\); default_zero(\$v6483\); 
          default_zero(\$12296\); default_zero(\$v3740\); 
          default_zero(\$11486\); default_zero(\$12040\); 
          default_zero(\$13252_c\); default_zero(\$v4919\); 
          default_zero(\$12292\); default_zero(\$10833\); 
          default_zero(\$v5772\); default_zero(\$v5165\); 
          default_zero(\$11821\); default_zero(\$v3872\); 
          default_zero(\$12893\); default_zero(\$v4228\); 
          default_zero(\$v5503\); default_zero(\$v5779\); 
          default_zero(\$v5628\); default_zero(\$v6432\); 
          default_zero(\$v4092\); default_zero(\$11848\); 
          default_zero(\$v5207\); default_zero(\$v4154\); 
          default_zero(\$v5970\); default_zero(\$13529_i\); 
          default_zero(\$v5480\); default_zero(\$v4152\); 
          default_zero(\$12042\); default_zero(\$v3838\); 
          default_zero(\$v4566\); default_zero(\$v3674\); 
          default_zero(\$14770\); default_zero(\$14404_i\); 
          default_zero(\$12876\); default_zero(\$v5240\); 
          default_zero(\$v6107\); default_zero(\$v6613\); 
          default_zero(\$v4291\); default_zero(\$15092\); 
          default_zero(\$v4840\); default_zero(\$v3374\); 
          default_zero(\$15479_i\); default_zero(\$v4625\); 
          default_zero(\$14795_i\); default_zero(\$v3806\); 
          default_zero(\$v6396\); default_zero(\$13086\); 
          default_zero(\$12030\); default_zero(\$v5981\); 
          default_zero(\$v4896\); default_zero(\$v3687\); 
          default_zero(\$v6592\); default_zero(\$v6010\); 
          default_zero(\$13808\); default_zero(\$v6380\); 
          default_zero(\$v6224\); default_zero(\$v5438\); 
          default_zero(\$v4244\); default_zero(\$15294\); 
          default_zero(\$v6349\); default_zero(\$13351\); 
          default_zero(\$11303\); default_zero(\$v5896\); 
          default_zero(\$v3936\); default_zero(\$v6957\); 
          default_zero(\$15636\); default_zero(\$13408\); 
          default_zero(\$10819\); default_zero(\$v3395\); 
          default_zero(\$12559\); default_zero(\$v6570\); 
          default_zero(\$v5861\); default_zero(\$12398_i\); 
          default_zero(\$v4685\); default_zero(\$v6408\); 
          default_zero(\$12610_j\); default_zero(\$v3388\); 
          default_zero(\$12311\); default_zero(\$v3900\); 
          default_zero(\$v4693\); default_zero(\$14533_opnd\); 
          default_zero(\$v6127\); default_zero(\$v3475\); 
          default_zero(\$v4020\); default_zero(\$v4961\); 
          default_zero(\$12248_i\); default_zero(\$v5643\); 
          default_zero(\$v4803\); default_zero(\$v5754\); 
          default_zero(\$11558\); default_zero(\$15263_i\); 
          default_zero(\$v4687\); default_zero(\$v5965\); 
          default_zero(\$v4966\); default_zero(\$12798\); 
          default_zero(\$14912\); default_zero(\$12177\); 
          default_zero(\$v3953\); default_zero(\$v4037\); 
          default_zero(\$v6821\); 
          default_zero(\$14863_list_tail2653331_arg\); 
          default_zero(\$v4509\); default_zero(\$v4046\); 
          default_zero(\$v5953\); default_zero(\$v3705\); 
          default_zero(\$12608_i\); default_zero(\$v3431\); 
          default_zero(\$14248\); default_zero(\$v6575\); 
          default_zero(\$12185\); default_zero(\$v4281\); 
          default_zero(\$v6019\); default_zero(\$14892_i\); 
          default_zero(\$12186\); default_zero(\$v4637\); 
          default_zero(\$15454\); default_zero(\$v4804\); 
          default_zero(\$11560_i\); default_zero(\$v5323\); 
          default_zero(\$v4515\); default_zero(\$v4340\); 
          default_zero(\$v6139\); default_zero(\$11482_i\); 
          default_zero(\$v6384\); default_zero(\$v5892\); 
          default_zero(\$v3932\); default_zero(\$v6625\); 
          default_zero(\$14720_i\); default_zero(\$11814\); 
          default_zero(\$v5509\); default_zero(\$11042\); 
          default_zero(\$v4830\); default_zero(\$13607\); 
          default_zero(\$v3486\); default_zero(\$v4511\); 
          default_zero(\$v4329\); default_zero(\$v3889\); 
          default_zero(\$15032\); default_zero(\$v6336\); 
          default_zero(\$v3719\); default_zero(\$15673\); 
          default_zero(\$v4900\); default_zero(\$v6309\); 
          default_zero(\$12471_i\); default_zero(\$v5586\); 
          default_zero(\$12297_x\); default_zero(\$13600_i\); 
          default_zero(\$13718_i\); default_zero(\$v3681\); 
          default_zero(\$v5776\); default_zero(\$v6469\); 
          default_zero(\$v6351\); default_zero(\$v4033\); 
          default_zero(\$15186_i\); default_zero(\$14719_i\); 
          default_zero(\$v5515\); default_zero(\$v3748\); 
          default_zero(\$v6404\); default_zero(\$v4769\); 
          default_zero(\$14772\); default_zero(\$12888\); 
          default_zero(\$13999_i\); default_zero(\$v4058\); 
          default_zero(\$v5363\); default_zero(\$v5632\); 
          default_zero(\$v4218\); default_zero(\$v4979\); 
          default_zero(\$11812\); default_zero(\$v6572\); 
          default_zero(\$v6376\); default_zero(\$11148\); 
          default_zero(\$v5119\); default_zero(\$v6652\); 
          default_zero(\$v6372\); default_zero(\$11748_i\); 
          default_zero(\$12786\); default_zero(\$v4853\); 
          default_zero(\$v4265\); default_zero(\$v6273\); 
          default_zero(\$v5764\); default_zero(\$13640_i\); 
          default_zero(\$v4611\); default_zero(\$15640\); 
          default_zero(\$v4727\); default_zero(\$v6091\); 
          default_zero(\$15555_len_aux3143354_result\); 
          default_zero(\$v3596\); default_zero(\$v4205\); 
          default_zero(\$v5828\); default_zero(\$v4481\); 
          default_zero(\$13546\); default_zero(\$v4728\); 
          default_zero(\$v4596\); default_zero(\$v3411\); 
          default_zero(\$14603\); default_zero(\$13405\); 
          default_zero(\$v6560\); default_zero(\$v4287\); 
          default_zero(\$v4845\); default_zero(\$v3965\); 
          default_zero(\$13744\); default_zero(\$v3547\); 
          default_zero(\$11449\); default_zero(\$v5058\); 
          default_zero(\$13222\); default_zero(\$v6936\); 
          default_zero(\$10740\); default_zero(\$v5052\); 
          default_zero(\$15702\); default_zero(\$15141\); 
          default_zero(\$15034_i\); default_zero(\$11121_i\); 
          default_zero(\$14650\); default_zero(\$13972\); 
          default_zero(\$v3910\); default_zero(\$v4936\); 
          default_zero(\$15293\); default_zero(\$v5413\); 
          default_zero(\$v4579\); default_zero(\$v6298\); 
          default_zero(\$v5702\); default_zero(\$12755_i\); 
          default_zero(\$v3682\); default_zero(\$v5481\); 
          default_zero(\$v5609\); default_zero(\$v5288\); 
          default_zero(\$12828_b\); default_zero(\$10749\); 
          default_zero(\$13606\); default_zero(\$v5261\); 
          default_zero(\$12348_i\); default_zero(\$v6664\); 
          default_zero(\$v3633\); default_zero(\$v5331\); 
          default_zero(\$v6633\); default_zero(\$v3637\); 
          default_zero(\$v4695\); default_zero(\$v4888\); 
          default_zero(\$v6235\); default_zero(\$12955_i\); 
          default_zero(\$v5348\); default_zero(\$13415\); 
          default_zero(\$v3429\); default_zero(\$14072_i\); 
          default_zero(\$v4908\); default_zero(\$v6668\); 
          default_zero(\$12685\); default_zero(\$v5120\); 
          default_zero(\$v3503\); 
          default_zero(\$13318_list_tail2653256_arg\); 
          default_zero(\$13178_i\); default_zero(\$v4988\); 
          default_zero(\$v5388\); default_zero(\$v4680\); 
          default_zero(\$14017\); default_zero(\$13667\); 
          default_zero(\$11571\); default_zero(result3365); 
          default_zero(\$v4691\); default_zero(\$v4745\); 
          default_zero(\$v3483\); default_zero(\$11903_i\); 
          default_zero(\$v6737\); default_zero(\$v4805\); 
          default_zero(\$v5823\); default_zero(\$15314\); 
          default_zero(\$14839\); default_zero(\$15071\); 
          default_zero(\$v5831\); default_zero(\$13155_i\); 
          default_zero(\$v6161\); default_zero(\$v4595\); 
          default_zero(\$v5308\); default_zero(\$v4601\); 
          default_zero(\$v6838\); default_zero(\$v6621\); 
          default_zero(\$15788_get_int268_result\); default_zero(\$v6108\); 
          default_zero(\$v5321\); default_zero(\$v4817\); 
          default_zero(\$v6392\); default_zero(\$v6304\); 
          default_zero(\$v6916\); default_zero(\$v4236\); 
          default_zero(\$v4878\); default_zero(\$v6739\); 
          default_zero(\$13461\); default_zero(\$v5380\); 
          default_zero(\$v5392\); default_zero(\$13596_v\); 
          default_zero(\$v6676\); default_zero(\$v3592\); 
          default_zero(\$v3653\); default_zero(\$11214\); 
          default_zero(\$v3456\); default_zero(\$11006_i\); 
          default_zero(\$11196_loop2913158_arg\); default_zero(\$v6492\); 
          default_zero(\$12880\); default_zero(\$14858_i\); 
          default_zero(\$v4197\); default_zero(\$15217_loop1312_arg\); 
          default_zero(\$v6413\); default_zero(\$11756\); 
          default_zero(\$11065_i\); default_zero(\$v7018\); 
          default_zero(\$10980\); default_zero(\$v5382\); 
          default_zero(\$12990_i\); default_zero(\$v5157\); 
          default_zero(\$v5943\); default_zero(\$13295\); 
          default_zero(\$v5124\); default_zero(\$v4623\); 
          default_zero(\$v6710\); default_zero(\$15033\); 
          default_zero(\$v3621\); default_zero(\$v5370\); 
          default_zero(\$v3660\); default_zero(\$12494_i\); 
          default_zero(\$10793\); default_zero(\$12790_i\); 
          default_zero(\$11803\); default_zero(\$10731\); 
          default_zero(\$v5771\); default_zero(\$v6555\); 
          default_zero(\$v5223\); default_zero(\$v6254\); 
          default_zero(\$13129_a\); default_zero(\$v5856\); 
          default_zero(\$11236\); default_zero(\$13741\); 
          default_zero(\$v3499\); default_zero(\$v3416\); 
          default_zero(\$v5810\); 
          default_zero(\$15724_len_aux3143361_result\); 
          default_zero(\$v3991\); default_zero(\$v4469\); 
          default_zero(\$v6303\); default_zero(\$11172_i\); 
          default_zero(\$12598\); default_zero(\$12556_i\); 
          default_zero(\$v3375\); default_zero(\$v6706\); 
          default_zero(\$v3893\); default_zero(\$v4967\); 
          default_zero(\$v5173\); default_zero(\$12105\); 
          default_zero(\$14834_i\); default_zero(\$15755\); 
          default_zero(\$11327\); default_zero(\$v5130\); 
          default_zero(\$v5954\); default_zero(\$v3539\); 
          default_zero(\$v6803\); default_zero(\$v6203\); 
          default_zero(\$10842\); default_zero(\$11333\); 
          default_zero(\$v4364\); default_zero(\$v4729\); 
          default_zero(\$v4210\); default_zero(\$v4588\); 
          default_zero(\$v3894\); default_zero(\$v5397\); 
          default_zero(\$v4308\); default_zero(\$15137\); 
          default_zero(\$12788\); default_zero(\$v6445\); 
          default_zero(\$15240_loop23133355_arg\); default_zero(\$14540\); 
          default_zero(\$v3600\); default_zero(\$14974\); 
          default_zero(\$v5269\); default_zero(\$v3836\); 
          default_zero(\$v6246\); default_zero(\$v5324\); 
          default_zero(\$12928_b\); default_zero(\$v4355\); 
          default_zero(\$v6117\); default_zero(\$v6825\); 
          default_zero(\$v5317\); default_zero(\$v3551\); 
          default_zero(\$11328_cont\); default_zero(\$v3514\); 
          default_zero(\$v4473\); default_zero(\$v6261\); 
          default_zero(\$12031\); default_zero(\$v4688\); 
          default_zero(\$12545\); default_zero(\$v5346\); 
          default_zero(\$v3752\); default_zero(\$13868_j\); 
          default_zero(\$v5043\); default_zero(\$12597\); 
          default_zero(\$v6681\); default_zero(\$12041_i\); 
          default_zero(\$10981\); default_zero(\$v4415\); 
          default_zero(\$14558\); default_zero(\$14705_i\); 
          default_zero(\$v6609\); default_zero(\$v3500\); 
          default_zero(\$v6112\); default_zero(\$v4726\); 
          default_zero(\$v4944\); default_zero(\$v5125\); 
          default_zero(\$12313\); default_zero(\$v4645\); 
          default_zero(\$v5329\); default_zero(\$v6794\); 
          default_zero(\$14284_i\); default_zero(\$15733\); 
          default_zero(\$11520_i\); default_zero(\$v4570\); 
          default_zero(\$v5778\); default_zero(\$10726\); 
          default_zero(\$13750\); default_zero(\$v4724\); 
          default_zero(\$v6255\); 
          default_zero(\$14863_list_tail2653331_result\); 
          default_zero(\$11966\); default_zero(\$15629\); 
          default_zero(\$v6269\); default_zero(\$15471_i\); 
          default_zero(\$14458_i\); default_zero(\$v3992\); 
          default_zero(\$v4669\); default_zero(\$v5568\); 
          default_zero(\$15324\); default_zero(\$v5496\); 
          default_zero(\$v6252\); default_zero(\$15506\); 
          default_zero(\$v3422\); default_zero(\$v5349\); 
          default_zero(\$14158_i\); default_zero(\$12993\); 
          default_zero(\$v6165\); default_zero(\$v6182\); 
          default_zero(\$v5618\); default_zero(\$12309\); 
          default_zero(\$v3490\); default_zero(\$v5354\); 
          default_zero(\$v3383\); default_zero(\$v6782\); 
          default_zero(\$v6364\); default_zero(\$v3860\); 
          default_zero(\$v6605\); default_zero(\$v4701\); 
          default_zero(\$v4495\); default_zero(\$v5147\); 
          default_zero(\$12299\); default_zero(\$v3980\); 
          default_zero(\$v5730\); default_zero(\$v5007\); 
          default_zero(\$v6116\); default_zero(\$v5570\); 
          default_zero(\$v4777\); default_zero(\$12300\); 
          default_zero(\$v3430\); default_zero(\$14390_i\); 
          default_zero(\$v5047\); default_zero(\$v3915\); 
          default_zero(\$v5294\); default_zero(\$15240_loop23133355_result\); 
          default_zero(\$13509\); default_zero(\$v5266\); 
          default_zero(\$15431_i\); default_zero(\$v5189\); 
          default_zero(\$14643\); default_zero(\$12855_i\); 
          default_zero(\$12113\); default_zero(\$13985_i\); 
          default_zero(\$12473\); default_zero(\$10897_k\); 
          default_zero(\$v5780\); default_zero(\$v5809\); 
          default_zero(\$v3387\); default_zero(\$v4090\); 
          default_zero(\$12614_i\); default_zero(\$10814\); 
          default_zero(\$13128_b\); default_zero(\$v6569\); 
          default_zero(\$v6590\); default_zero(\$14185_i\); 
          default_zero(\$11321_i\); default_zero(\$11730\); 
          default_zero(\$12985_y\); default_zero(\$v5747\); 
          default_zero(\$v4609\); default_zero(\$v5468\); 
          default_zero(\$v4402\); default_zero(\$14763_i\); 
          default_zero(\$12414\); default_zero(\$v6400\); 
          default_zero(\$v6388\); default_zero(\$v3577\); 
          default_zero(\$15763_j\); default_zero(\$11962\); 
          default_zero(\$v6478\); default_zero(\$15068_opnd\); 
          default_zero(\$v6961\); default_zero(\$v6998\); 
          default_zero(\$v5169\); default_zero(\$v6979\); 
          default_zero(\$v5090\); default_zero(\$v3689\); 
          default_zero(\$v3543\); 
          default_zero(\$14481_decode_loop310_result\); 
          default_zero(\$v3701\); default_zero(\$v5523\); 
          default_zero(\$14580_i\); default_zero(\$v4180\); 
          default_zero(\$v3535\); default_zero(\$13829_i\); 
          default_zero(\$12420_x\); default_zero(\$v5098\); 
          default_zero(\$v6809\); default_zero(\$v4438\); 
          default_zero(\$v5873\); default_zero(\$15465\); 
          default_zero(\$v4147\); default_zero(\$12104\); 
          default_zero(\$v3373\); default_zero(\$v5390\); 
          default_zero(\$v4885\); default_zero(\$v6579\); 
          default_zero(\$12785_y\); default_zero(\$14080\); 
          default_zero(\$v5053\); default_zero(\$v3465\); 
          default_zero(\$11147_i\); default_zero(\$v6584\); 
          default_zero(\$v6289\); default_zero(\$v6066\); 
          default_zero(\$14409\); default_zero(\$v5482\); 
          default_zero(\$v4424\); default_zero(\$14972\); 
          default_zero(\$v5959\); default_zero(\$15261\); 
          default_zero(\$13832\); default_zero(\$v3448\); 
          default_zero(\$v5077\); default_zero(\$v6912\); 
          default_zero(\$12433_i\); default_zero(\$12083_i\); 
          default_zero(\$15129_i\); default_zero(\$10900\); 
          default_zero(\$14722\); default_zero(\$v6817\); 
          default_zero(\$15303_str_rib\); default_zero(\$v6799\); 
          default_zero(\$v6994\); default_zero(\$15091\); 
          default_zero(\$v4346\); default_zero(\$v6424\); 
          default_zero(\$v6421\); default_zero(\$15555_len_aux3143354_arg\); 
          default_zero(\$12431\); default_zero(\$10721\); 
          default_zero(\$v4554\); default_zero(\$v6525\); 
          default_zero(\$v5036\); default_zero(\$v5121\); 
          default_zero(\$v3678\); default_zero(\$14079\); 
          default_zero(\$v6245\); default_zero(\$v5011\); 
          default_zero(\$v6918\); default_zero(\$v4546\); 
          default_zero(\$13291_i\); default_zero(\$v4915\); 
          default_zero(\$14662\); default_zero(\$v4086\); 
          default_zero(\$v4042\); default_zero(\$12169\); 
          default_zero(\$14306\); default_zero(\$13234\); 
          default_zero(\$v3565\); default_zero(\$v5799\); 
          default_zero(\$v6846\); default_zero(\$11655_i\); 
          default_zero(\$v6863\); default_zero(\$v5289\); 
          default_zero(\$12976\); default_zero(\$11787_i\); 
          default_zero(\$11437_loop3073170_arg\); default_zero(\$v6897\); 
          default_zero(\$13626_i\); default_zero(\$v4653\); 
          default_zero(\$v4260\); default_zero(\$12980\); 
          default_zero(\$v3661\); default_zero(\$11665\); 
          default_zero(\$10979_i\); default_zero(\$v4678\); 
          default_zero(\$13177\); default_zero(\$11658\); 
          default_zero(\$12972\); default_zero(\$15796\); 
          default_zero(\$15613_i\); default_zero(\$v3896\); 
          default_zero(\$11406_i\); default_zero(\$v4360\); 
          default_zero(\$v6646\); default_zero(\$v5365\); 
          default_zero(\$v4380\); default_zero(\$v3928\); 
          default_zero(\$v3381\); default_zero(\$v4679\); 
          default_zero(\$12261_i\); default_zero(\$14897_get_int268_arg\); 
          default_zero(\$10766\); default_zero(\$v4957\); 
          default_zero(\$v6965\); default_zero(\$v5040\); 
          default_zero(\$12879\); default_zero(\$15788_get_int268_arg\); 
          default_zero(\$v6940\); default_zero(\$v3717\); 
          default_zero(\$v5872\); default_zero(\$v4712\); 
          default_zero(\$13296\); default_zero(\$v4502\); 
          default_zero(\$v4802\); default_zero(\$v6766\); 
          default_zero(\$v5633\); default_zero(\$14658\); 
          default_zero(\$v4973\); default_zero(\$v6122\); 
          default_zero(\$v3463\); default_zero(\$v3376\); 
          default_zero(\$12587\); default_zero(\$14681_i\); 
          default_zero(\$v5552\); default_zero(\$v4589\); 
          default_zero(\$v6535\); default_zero(\$v6660\); 
          default_zero(\$14648_ty\); default_zero(\$11713\); 
          default_zero(\$v6922\); default_zero(\$v5696\); 
          default_zero(\$12543_x\); default_zero(\$v3567\); 
          default_zero(\$v3736\); default_zero(\$12678_x\); 
          default_zero(\$v5822\); default_zero(\$v4861\); 
          default_zero(\$v6718\); default_zero(\$v3417\); 
          default_zero(\$v3715\); default_zero(\$v5198\); 
          default_zero(\$v4172\); default_zero(\$v3773\); 
          default_zero(\$v5837\); default_zero(\$v6441\); 
          default_zero(\$11596\); default_zero(\$v5563\); 
          default_zero(\$11905\); default_zero(\$v5337\); 
          default_zero(\$14211_i\); default_zero(\$v4684\); 
          default_zero(\$14683\); default_zero(\$12110_i\); 
          default_zero(\$v4141\); default_zero(\$14595_i\); 
          default_zero(\$v5073\); default_zero(\$v6521\); 
          default_zero(\$v6033\); default_zero(\$v3753\); 
          default_zero(\$13482_i\); default_zero(\$v3531\); 
          default_zero(\$12035\); default_zero(\$15611_i\); 
          default_zero(\$v4709\); default_zero(\$v5492\); 
          default_zero(\$v3843\); default_zero(\$14837\); 
          default_zero(\$12415\); default_zero(\$v4155\); 
          default_zero(\$v6901\); default_zero(\$v5727\); 
          default_zero(\$v5463\); default_zero(\$14415\); 
          default_zero(\$v3527\); default_zero(\$v4602\); 
          default_zero(\$15313\); default_zero(\$v5725\); 
          default_zero(\$v4750\); default_zero(\$v3667\); 
          default_zero(\$v5068\); default_zero(\$12305_y\); 
          default_zero(\$v4101\); default_zero(\$v4465\); 
          default_zero(\$11433_i\); default_zero(\$v6352\); 
          default_zero(\$11213\); default_zero(\$15298\); 
          default_zero(rdy3363); default_zero(\$12190\); 
          default_zero(\$12225_i\); default_zero(\$11280_i\); 
          default_zero(\$v5133\); default_zero(\$v5734\); 
          default_zero(\$12607_j\); default_zero(\$v3769\); 
          default_zero(\$v4025\); default_zero(\$10828_c2_rib\); 
          default_zero(\$v5832\); default_zero(\$v3793\); 
          default_zero(\$10767_j\); default_zero(\$15306\); 
          default_zero(\$v4347\); default_zero(\$v6893\); 
          default_zero(\$15760_i\); default_zero(\$12053\); 
          default_zero(\$v6714\); default_zero(\$v6325\); 
          default_zero(\$14936\); default_zero(\$v6236\); 
          default_zero(\$v6330\); default_zero(\$v4994\); 
          default_zero(\$11675\); default_zero(\$v6449\); 
          default_zero(\$10750\); default_zero(\$v5275\); 
          default_zero(\$13085_y\); default_zero(\$v5830\); 
          default_zero(\$v4339\); default_zero(\$v5975\); 
          default_zero(\$v5260\); default_zero(\$v4532\); 
          default_zero(\$v5726\); default_zero(\$v5976\); 
          default_zero(\$v4825\); default_zero(\$13665\); 
          default_zero(\$15467_str_rib\); default_zero(\$v4558\); 
          default_zero(\$14301\); default_zero(\$v5259\); 
          default_zero(\$v5141\); default_zero(\$v4681\); 
          default_zero(\$v5748\); default_zero(\$11543\); 
          default_zero(\$11972_i\); default_zero(\$v3940\); 
          default_zero(\$v4449\); default_zero(\$v6359\); 
          default_zero(\$v7010\); default_zero(\$12122\); 
          default_zero(\$v5335\); default_zero(\$v4217\); 
          default_zero(\$v4388\); default_zero(\$11971\); 
          default_zero(\$v4457\); default_zero(\$v6795\); 
          default_zero(\$11736_x\); default_zero(\$14472_i\); 
          default_zero(\$v5560\); default_zero(\$v4932\); 
          default_zero(\$v4751\); default_zero(\$v4911\); 
          default_zero(\$v6875\); default_zero(\$10893_i\); 
          default_zero(\$13028_b\); default_zero(\$v5508\); 
          default_zero(\$14541\); default_zero(\$v3578\); 
          default_zero(\$v5597\); default_zero(\$v6072\); 
          default_zero(\$v6073\); default_zero(\$v4718\); 
          default_zero(\$v5102\); default_zero(\$v5694\); 
          default_zero(\$v6578\); default_zero(\$v3552\); 
          default_zero(\$v3447\); default_zero(\$11134_i\); 
          default_zero(\$15457\); default_zero(\$11548_y\); 
          default_zero(\$v6859\); default_zero(\$12889\); 
          default_zero(\$v6216\); default_zero(\$v4990\); 
          default_zero(\$v3580\); default_zero(\$v6689\); 
          default_zero(\$v4000\); default_zero(\$15262\); 
          default_zero(\$v5502\); default_zero(\$v5276\); 
          default_zero(\$14840\); default_zero(\$13869_i\); 
          default_zero(\$14405_i\); default_zero(\$12984\); 
          default_zero(\$11809\); default_zero(\$v6305\); 
          default_zero(\$11047\); default_zero(\$13837\); 
          default_zero(\$v4702\); default_zero(\$v3716\); 
          default_zero(\$v6135\); default_zero(\$v4016\); 
          default_zero(\$13967\); default_zero(\$11819\); 
          default_zero(\$v4168\); default_zero(\$v3848\); 
          default_zero(\$v3924\); default_zero(\$v5356\); 
          default_zero(\$v5391\); default_zero(\$v3585\); 
          default_zero(\$15319\); default_zero(\$v5821\); 
          default_zero(\$v4810\); default_zero(\$v4270\); 
          default_zero(\$11667_i\); default_zero(\$v3672\); 
          default_zero(\$11738\); default_zero(\$v7014\); 
          default_zero(\$13595_i\); default_zero(\$v6685\); 
          default_zero(\$11657\); default_zero(\$v6580\); 
          default_zero(\$15475_end_rib\); default_zero(\$v4252\); 
          default_zero(\$10765\); default_zero(\$12776\); 
          default_zero(\$v4085\); default_zero(\$v5146\); 
          default_zero(\$v4698\); default_zero(\$13872_j\); 
          default_zero(\$12670_i\); default_zero(\$v3484\); 
          default_zero(\$v6754\); default_zero(\$12616_j\); 
          default_zero(\$11708\); default_zero(\$v3807\); 
          default_zero(\$v4422\); default_zero(\$v5709\); 
          default_zero(\$v5231\); default_zero(\$v3469\); 
          default_zero(\$v3493\); default_zero(\$v4608\); 
          default_zero(\$v4423\); default_zero(\$v4550\); 
          default_zero(\$v4794\); default_zero(\$15473\); 
          default_zero(\$v4128\); default_zero(\$14872\); 
          default_zero(\$v3504\); default_zero(\$v5548\); 
          default_zero(\$v3808\); default_zero(\$v3458\); 
          default_zero(\$15598_j\); default_zero(\$v5336\); 
          default_zero(\$12599_i\); default_zero(\$v4398\); 
          default_zero(\$v4983\); default_zero(\$15434_j\); 
          default_zero(\$v3400\); default_zero(\$13545_i\); 
          default_zero(\$v5156\); default_zero(\$v5454\); 
          default_zero(\$v6526\); default_zero(\$15564\); 
          default_zero(\$v6285\); default_zero(\$12691_i\); 
          default_zero(\$v6099\); default_zero(\$v3732\); 
          default_zero(\$v4403\); default_zero(\$11448\); 
          default_zero(\$11228_i\); default_zero(\$11293_i\); 
          default_zero(\$v6045\); default_zero(\$v4836\); 
          default_zero(\$v6140\); default_zero(\$11551\); 
          default_zero(\$v4216\); default_zero(\$v4694\); 
          default_zero(\$v5396\); default_zero(\$v5579\); 
          default_zero(\$15630_i\); default_zero(\$v4953\); 
          default_zero(\$v5353\); default_zero(\$13598\); 
          default_zero(\$v5051\); default_zero(\$v3724\); 
          default_zero(\$v6990\); default_zero(\$13460\); 
          default_zero(\$10737\); default_zero(\$11627_i\); 
          default_zero(\$12384_i\); default_zero(\$v6187\); 
          default_zero(\$v5720\); default_zero(\$v5556\); 
          default_zero(\$11944_i\); default_zero(\$12605_i\); 
          default_zero(\$v4857\); default_zero(\$v6756\); 
          default_zero(\$v6604\); default_zero(\$v5421\); 
          default_zero(\$15342\); default_zero(\$12173\); 
          default_zero(\$12971\); default_zero(\$15563\); 
          default_zero(\$15488\); default_zero(\$v4884\); 
          default_zero(\$v6332\); default_zero(\$11666\); 
          default_zero(\$14445_i\); default_zero(\$v3813\); 
          default_zero(\$v3457\); default_zero(\$v5791\); 
          default_zero(\$v3477\); default_zero(\$v6054\); 
          default_zero(\$v3636\); default_zero(\$14642\); 
          default_zero(\$11594\); default_zero(\$v3491\); 
          default_zero(\$v5569\); default_zero(\$v3972\); 
          default_zero(\$v5983\); default_zero(\$v6735\); 
          default_zero(\$v5126\); default_zero(\$12308\); 
          default_zero(\$v6315\); default_zero(\$v5881\); 
          default_zero(\$10848\); default_zero(\$v5827\); 
          default_zero(\$15131\); default_zero(\$v5387\); 
          default_zero(\$v6212\); default_zero(\$v4665\); 
          default_zero(\$v6638\); 
          default_zero(\$15391_len_aux3143348_result\); 
          default_zero(\$v3852\); default_zero(\$v3744\); 
          default_zero(\$v5190\); default_zero(\$12176\); 
          default_zero(\$12793\); default_zero(\$14939_get_int268_arg\); 
          default_zero(\$11670\); default_zero(\$v5495\); 
          default_zero(\$v5274\); default_zero(\$13684_i\); 
          default_zero(\$v5475\); default_zero(\$15628\); 
          default_zero(\$11668\); default_zero(\$11149\); 
          default_zero(\$v5561\); default_zero(\$11466_i\); 
          default_zero(\$11223\); default_zero(\$13216\); 
          default_zero(\$15734\); default_zero(\$12291\); 
          default_zero(\$v5982\); default_zero(\$v4630\); 
          default_zero(\$v3703\); default_zero(\$v6457\); 
          default_zero(\$11267_i\); default_zero(\$v4720\); 
          default_zero(\$v6577\); default_zero(\$15594_j\); 
          default_zero(\$v5562\); default_zero(\$v6377\); 
          default_zero(\$v5045\); default_zero(\$v4670\); 
          default_zero(\$14728\); default_zero(\$v5880\); 
          default_zero(\$13382_i\); default_zero(\$13769_i\); 
          default_zero(\$11709\); default_zero(\$v3455\); 
          default_zero(\$14651\); default_zero(\$12991\); 
          default_zero(\$v4137\); default_zero(\$v3470\); 
          default_zero(\$12304\); default_zero(\$12226\); 
          default_zero(\$v5341\); default_zero(\$15470\); 
          default_zero(\$13098\); default_zero(\$v4889\); 
          default_zero(\$v6368\); default_zero(\$v6231\); 
          default_zero(\$v5829\); default_zero(\$v5111\); 
          default_zero(\$v4256\); default_zero(\$v3643\); 
          default_zero(\$v6672\); default_zero(\$v5510\); 
          default_zero(\$v5848\); default_zero(\$13443_i\); 
          default_zero(\$v6422\); default_zero(\$v4372\); 
          default_zero(\$11504_i\); default_zero(\$v5701\); 
          default_zero(\$v5922\); default_zero(\$v5591\); 
          default_zero(\$v5531\); default_zero(\$v4600\); 
          default_zero(\$11826\); default_zero(\$v4626\); 
          default_zero(\$11380\); default_zero(\$v3659\); 
          default_zero(\$11048\); default_zero(\$v3412\); 
          default_zero(\$v5483\); default_zero(\$v6980\); 
          default_zero(\$13666\); default_zero(\$14192\); 
          default_zero(\$v5989\); default_zero(\$11218\); 
          default_zero(\$v5803\); default_zero(\$v6904\); 
          default_zero(\$v3709\); default_zero(\$v4883\); 
          default_zero(\$12686_y\); default_zero(\$v4583\); 
          default_zero(\$v4737\); default_zero(\$v6345\); 
          default_zero(\$v6571\); default_zero(\$v5268\); 
          default_zero(\$v6079\); default_zero(\$v5500\); 
          default_zero(\$v3683\); default_zero(\$14666\); 
          default_zero(\$12877_x\); default_zero(\$11219\); 
          default_zero(\$v4108\); default_zero(\$12604_j\); 
          default_zero(\$12428_y\); default_zero(\$v6123\); 
          default_zero(\$v5713\); default_zero(\$v5110\); 
          default_zero(\$v4526\); default_zero(\$v6833\); 
          default_zero(\$v6290\); default_zero(\$v3981\); 
          default_zero(\$v5871\); default_zero(\$v6573\); 
          default_zero(\$v3510\); default_zero(\$v4831\); 
          default_zero(\$11032_i\); default_zero(\$11535\); 
          default_zero(\$11420_i\); default_zero(\$14655\); 
          default_zero(\$13399\); default_zero(\$12039\); 
          default_zero(\$13327\); default_zero(\$14012_i\); 
          default_zero(\$v4024\); default_zero(\$10839_s\); 
          default_zero(\$v6807\); default_zero(\$v3647\); 
          default_zero(\$v5805\); default_zero(\$v6576\); 
          default_zero(\$v5403\); default_zero(\$v5297\); 
          default_zero(\$v3591\); default_zero(\$v6647\); 
          default_zero(\$11556_z\); default_zero(\$v5473\); 
          default_zero(\$v4987\); default_zero(\$v5887\); 
          default_zero(\$v6032\); default_zero(\$v3983\); 
          default_zero(\$v3497\); default_zero(\$13089\); 
          default_zero(\$12552\); default_zero(\$v6157\); 
          default_zero(\$11912\); default_zero(\$v5106\); 
          default_zero(\$13783_i\); default_zero(\$v6170\); 
          default_zero(\$v5242\); default_zero(\$v5381\); 
          default_zero(\$v4789\); default_zero(\$v5474\); 
          default_zero(\$v5062\); default_zero(\$11804\); 
          default_zero(\$v6153\); default_zero(\$v5718\); 
          default_zero(\$v4269\); default_zero(\$v3895\); 
          default_zero(\$v5906\); default_zero(\$11911\); 
          default_zero(\$15217_loop1312_result\); default_zero(\$v5939\); 
          default_zero(\$v5758\); default_zero(\$14271_i\); 
          default_zero(\$14511_loop311_result\); default_zero(\$v5882\); 
          default_zero(\$v6966\); default_zero(\$10792\); 
          default_zero(\$10913_i\); default_zero(\$v4989\); 
          default_zero(\$v5219\); default_zero(\$11437_loop3073170_result\); 
          default_zero(\$v6412\); default_zero(\$v5375\); 
          default_zero(\$v5898\); default_zero(\$v3966\); 
          default_zero(\$v5581\); default_zero(\$v5797\); 
          default_zero(\$v6915\); default_zero(\$11100\); 
          default_zero(\$14125_i\); default_zero(\$v5115\); 
          default_zero(\$v4657\); default_zero(\$14542_new_rib\); 
          default_zero(\$v6074\); default_zero(\$v5501\); 
          default_zero(\$v6248\); default_zero(\$v5236\); 
          default_zero(\$v3655\); default_zero(\$12872\); 
          default_zero(\$11576\); default_zero(\$v4706\); 
          default_zero(\$v4717\); default_zero(\$v3952\); 
          default_zero(\$v5728\); default_zero(\$v6191\); 
          default_zero(\$v6975\); default_zero(\$v5984\); 
          default_zero(\$v6564\); default_zero(\$v4283\); 
          default_zero(\$v3516\); default_zero(\$v5672\); 
          default_zero(\$10896\); default_zero(\$13225\); 
          default_zero(\$11534\); default_zero(\$v3409\); 
          default_zero(\$v4261\); default_zero(\$15678\); 
          default_zero(\$15595_i\); default_zero(\$13746\); 
          default_zero(\$12550\); default_zero(\$v4091\); 
          default_zero(\$v5676\); default_zero(\$10826\); 
          default_zero(\$v7002\); default_zero(\$v6745\); 
          default_zero(\$v5241\); default_zero(\$11222\); 
          default_zero(\$15076_new_rib\); default_zero(\$v5660\); 
          default_zero(\$v6952\); default_zero(\$13547\); 
          default_zero(\$v5877\); default_zero(\$v5680\); 
          default_zero(\$15644\); default_zero(\$v4575\); 
          default_zero(\$v6064\); default_zero(\$v4444\); 
          default_zero(\$v4477\); default_zero(\$v6634\); 
          default_zero(\$v4012\); default_zero(\$v4962\); 
          default_zero(\$v5681\); default_zero(\$v6903\); 
          default_zero(\$12989\); default_zero(\$v5910\); 
          default_zero(\$v4080\); default_zero(\$v4296\); 
          default_zero(\$v5902\); default_zero(\$v4212\); 
          default_zero(\$14058_i\); default_zero(\$12436\); 
          default_zero(\$15477\); default_zero(\$v3817\); 
          default_zero(\$10757\); default_zero(\$v5583\); 
          default_zero(\$v5746\); default_zero(\$12718_a\); 
          default_zero(\$12829_a\); default_zero(\$v4008\); 
          default_zero(\$v6465\); default_zero(\$v3476\); 
          default_zero(\$v6141\); default_zero(\$v6145\); 
          default_zero(\$v3828\); default_zero(\$11338\); 
          default_zero(\$v3368\); default_zero(\$v6879\); 
          default_zero(\$v5668\); default_zero(\$13743_i\); 
          default_zero(\$15128_i\); default_zero(\$12884\); 
          default_zero(\$v4829\); default_zero(\$v5854\); 
          default_zero(\$11443\); default_zero(\$v6310\); 
          default_zero(\$12777_x\); default_zero(\$v5886\); 
          default_zero(\$v5914\); default_zero(\$v5798\); 
          default_zero(\$v4708\); default_zero(\$v4624\); 
          default_zero(\$15648\); default_zero(\$13850_i\); 
          default_zero(\$v3868\); default_zero(\$15074\); 
          default_zero(\$v6488\); default_zero(\$v5215\); 
          default_zero(\$v4153\); default_zero(\$v5787\); 
          default_zero(\$15035\); default_zero(\$11917\); 
          default_zero(\$10966_i\); default_zero(\$v5729\); 
          default_zero(\$v4439\); default_zero(\$v6226\); 
          default_zero(\$v6357\); default_zero(\$v4808\); 
          default_zero(\$v5399\); default_zero(\$11749\); 
          default_zero(\$v4508\); default_zero(\$11663\); 
          default_zero(\$15469\); default_zero(\$15632\); 
          default_zero(\$v5298\); default_zero(\$15043\); 
          default_zero(\$12555\); default_zero(\$14319_i\); 
          default_zero(\$v6867\); default_zero(\$v5588\); 
          default_zero(\$14536\); default_zero(\$13663_i\); 
          default_zero(\$10753\); default_zero(\$v6944\); 
          default_zero(\$v4397\); default_zero(\$v4705\); 
          default_zero(\$15090_i\); default_zero(\$13807\); 
          default_zero(\$v3502\); default_zero(\$v6063\); 
          default_zero(\$14407\); default_zero(\$v4869\); 
          default_zero(\$v5590\); default_zero(\$12289_i\); 
          default_zero(\$v5714\); default_zero(\$14198\); 
          default_zero(\$v6317\); default_zero(\$12690\); 
          default_zero(\$15268\); default_zero(\$v6932\); 
          default_zero(\$14682\); default_zero(\$13093\); 
          default_zero(\$v5330\); default_zero(\$13294\); 
          default_zero(\$v3864\); 
          default_zero(\$13500_list_tail2653266_result\); 
          default_zero(\$v6028\); default_zero(\$v5535\); 
          default_zero(\$v5946\); default_zero(\$v5078\); 
          default_zero(rdy3366); default_zero(\$11889_i\); 
          default_zero(\$14647\); default_zero(\$v5547\); 
          default_zero(\$12427\); default_zero(\$v3428\); 
          default_zero(\$v3432\); default_zero(\$v6311\); 
          rdy <= "1";
          rdy3363 := "0";
          state <= compute3364;
          state_var7021 <= compute3367;
          
        else if run = '1' then
          case state is
          when \$10694_forever290\ =>
            state <= \$10694_forever290\;
          when compute3364 =>
            rdy3363 := eclat_false;
            case state_var7021 is
            when \$10704_forever290\ =>
              state_var7021 <= \$10704_forever290\;
            when \$10778_run286\ =>
              \$v5622\ := \$$10700_pc_ptr_take\;
              if \$v5622\(0) = '1' then
                state_var7021 <= q_wait5621;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5619;
              end if;
            when \$10801_forever3163135\ =>
              state_var7021 <= \$10805_forever3163133\;
            when \$10805_forever3163133\ =>
              state_var7021 <= \$10805_forever3163133\;
            when \$10859_forever3163136\ =>
              state_var7021 <= \$10863_forever3163133\;
            when \$10863_forever3163133\ =>
              state_var7021 <= \$10863_forever3163133\;
            when \$10872_forever3163137\ =>
              state_var7021 <= \$10876_forever3163133\;
            when \$10876_forever3163133\ =>
              state_var7021 <= \$10876_forever3163133\;
            when \$10885_forever3163138\ =>
              state_var7021 <= \$10889_forever3163133\;
            when \$10889_forever3163133\ =>
              state_var7021 <= \$10889_forever3163133\;
            when \$10905_forever3163139\ =>
              state_var7021 <= \$10909_forever3163133\;
            when \$10909_forever3163133\ =>
              state_var7021 <= \$10909_forever3163133\;
            when \$10932_forever3163140\ =>
              state_var7021 <= \$10936_forever3163133\;
            when \$10936_forever3163133\ =>
              state_var7021 <= \$10936_forever3163133\;
            when \$10945_forever3163141\ =>
              state_var7021 <= \$10949_forever3163133\;
            when \$10949_forever3163133\ =>
              state_var7021 <= \$10949_forever3163133\;
            when \$10958_forever3163142\ =>
              state_var7021 <= \$10962_forever3163133\;
            when \$10962_forever3163133\ =>
              state_var7021 <= \$10962_forever3163133\;
            when \$10971_forever3163143\ =>
              state_var7021 <= \$10975_forever3163133\;
            when \$10975_forever3163133\ =>
              state_var7021 <= \$10975_forever3163133\;
            when \$10998_forever3163144\ =>
              state_var7021 <= \$11002_forever3163133\;
            when \$11002_forever3163133\ =>
              state_var7021 <= \$11002_forever3163133\;
            when \$11011_forever3163145\ =>
              state_var7021 <= \$11015_forever3163133\;
            when \$11015_forever3163133\ =>
              state_var7021 <= \$11015_forever3163133\;
            when \$11024_forever3163146\ =>
              state_var7021 <= \$11028_forever3163133\;
            when \$11028_forever3163133\ =>
              state_var7021 <= \$11028_forever3163133\;
            when \$11036_loop3073149\ =>
              \$v3509\ := \$11036_loop3073149_arg\(0 to 35);
              \$v3510\ := \$v3509\(0 to 3);
              \$v3504\ := \$v3509\(4 to 35);
              case \$v3510\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11073_forever3163148\;
              when "0000" =>
                \$11081_i\ := \$v3504\(0 to 31);
                \$v3508\ := \$$10696_ram_ptr_take\;
                if \$v3508\(0) = '1' then
                  state_var7021 <= q_wait3507;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11081_i\));
                  state_var7021 <= pause_getI3505;
                end if;
              when others =>
                
              end case;
            when \$11057_forever3163147\ =>
              state_var7021 <= \$11061_forever3163133\;
            when \$11061_forever3163133\ =>
              state_var7021 <= \$11061_forever3163133\;
            when \$11073_forever3163148\ =>
              state_var7021 <= \$11077_forever3163133\;
            when \$11077_forever3163133\ =>
              state_var7021 <= \$11077_forever3163133\;
            when \$11090_forever3163150\ =>
              state_var7021 <= \$11094_forever3163133\;
            when \$11094_forever3163133\ =>
              state_var7021 <= \$11094_forever3163133\;
            when \$11113_forever3163151\ =>
              state_var7021 <= \$11117_forever3163133\;
            when \$11117_forever3163133\ =>
              state_var7021 <= \$11117_forever3163133\;
            when \$11126_forever3163152\ =>
              state_var7021 <= \$11130_forever3163133\;
            when \$11130_forever3163133\ =>
              state_var7021 <= \$11130_forever3163133\;
            when \$11139_forever3163153\ =>
              state_var7021 <= \$11143_forever3163133\;
            when \$11143_forever3163133\ =>
              state_var7021 <= \$11143_forever3163133\;
            when \$11164_forever3163154\ =>
              state_var7021 <= \$11168_forever3163133\;
            when \$11168_forever3163133\ =>
              state_var7021 <= \$11168_forever3163133\;
            when \$11177_forever3163155\ =>
              state_var7021 <= \$11181_forever3163133\;
            when \$11181_forever3163133\ =>
              state_var7021 <= \$11181_forever3163133\;
            when \$11196_loop2913158\ =>
              \$v3576\ := eclat_eq(\$11196_loop2913158_arg\(0 to 31) & X"0000000" & X"0");
              if \$v3576\(0) = '1' then
                \$11196_loop2913158_result\ := \$11196_loop2913158_arg\(32 to 67);
                \$10839_s\ := \$11196_loop2913158_result\;
                \$v3517\ := \$10814\(72 to 107);
                \$v3518\ := \$v3517\(0 to 3);
                \$v3516\ := \$v3517\(4 to 35);
                case \$v3518\ is
                when "0001" =>
                  \$10840\ := eclat_false;
                when "0000" =>
                  \$11187_i\ := \$v3516\(0 to 31);
                  \$10840\ := eclat_if(eclat_ge(\$11187_i\ & X"0000000" & X"0") & eclat_lt(\$11187_i\ & X"0000" & X"2710") & eclat_false);
                when others =>
                  
                end case;
                \$v3515\ := \$10840\;
                if \$v3515\(0) = '1' then
                  \$v3436\ := \$$10697_stack_ptr_take\;
                  if \$v3436\(0) = '1' then
                    state_var7021 <= q_wait3435;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI3433;
                  end if;
                else
                  \$v3514\ := \$$10697_stack_ptr_take\;
                  if \$v3514\(0) = '1' then
                    state_var7021 <= q_wait3513;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI3511;
                  end if;
                end if;
              else
                \$v3575\ := \$$10697_stack_ptr_take\;
                if \$v3575\(0) = '1' then
                  state_var7021 <= q_wait3574;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3572;
                end if;
              end if;
            when \$11244_forever3163156\ =>
              state_var7021 <= \$11248_forever3163133\;
            when \$11248_forever3163133\ =>
              state_var7021 <= \$11248_forever3163133\;
            when \$11259_forever3163157\ =>
              state_var7021 <= \$11263_forever3163133\;
            when \$11263_forever3163133\ =>
              state_var7021 <= \$11263_forever3163133\;
            when \$11272_forever3163159\ =>
              state_var7021 <= \$11276_forever3163133\;
            when \$11276_forever3163133\ =>
              state_var7021 <= \$11276_forever3163133\;
            when \$11285_forever3163160\ =>
              state_var7021 <= \$11289_forever3163133\;
            when \$11289_forever3163133\ =>
              state_var7021 <= \$11289_forever3163133\;
            when \$11311_forever3163161\ =>
              state_var7021 <= \$11315_forever3163133\;
            when \$11315_forever3163133\ =>
              state_var7021 <= \$11315_forever3163133\;
            when \$11343_forever3163162\ =>
              state_var7021 <= \$11347_forever3163133\;
            when \$11347_forever3163133\ =>
              state_var7021 <= \$11347_forever3163133\;
            when \$11356_forever3163163\ =>
              state_var7021 <= \$11360_forever3163133\;
            when \$11360_forever3163133\ =>
              state_var7021 <= \$11360_forever3163133\;
            when \$11370_forever3163164\ =>
              state_var7021 <= \$11374_forever3163133\;
            when \$11374_forever3163133\ =>
              state_var7021 <= \$11374_forever3163133\;
            when \$11398_forever3163165\ =>
              state_var7021 <= \$11402_forever3163133\;
            when \$11402_forever3163133\ =>
              state_var7021 <= \$11402_forever3163133\;
            when \$11412_forever3163166\ =>
              state_var7021 <= \$11416_forever3163133\;
            when \$11416_forever3163133\ =>
              state_var7021 <= \$11416_forever3163133\;
            when \$11425_forever3163167\ =>
              state_var7021 <= \$11429_forever3163133\;
            when \$11429_forever3163133\ =>
              state_var7021 <= \$11429_forever3163133\;
            when \$11437_loop3073170\ =>
              \$v3710\ := \$11437_loop3073170_arg\(0 to 35);
              \$v3711\ := \$v3710\(0 to 3);
              \$v3705\ := \$v3710\(4 to 35);
              case \$v3711\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11474_forever3163169\;
              when "0000" =>
                \$11482_i\ := \$v3705\(0 to 31);
                \$v3709\ := \$$10696_ram_ptr_take\;
                if \$v3709\(0) = '1' then
                  state_var7021 <= q_wait3708;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11482_i\));
                  state_var7021 <= pause_getI3706;
                end if;
              when others =>
                
              end case;
            when \$11458_forever3163168\ =>
              state_var7021 <= \$11462_forever3163133\;
            when \$11462_forever3163133\ =>
              state_var7021 <= \$11462_forever3163133\;
            when \$11474_forever3163169\ =>
              state_var7021 <= \$11478_forever3163133\;
            when \$11478_forever3163133\ =>
              state_var7021 <= \$11478_forever3163133\;
            when \$11496_forever3163171\ =>
              state_var7021 <= \$11500_forever3163133\;
            when \$11500_forever3163133\ =>
              state_var7021 <= \$11500_forever3163133\;
            when \$11510_forever3163172\ =>
              state_var7021 <= \$11514_forever3163133\;
            when \$11514_forever3163133\ =>
              state_var7021 <= \$11514_forever3163133\;
            when \$11525_forever3163173\ =>
              state_var7021 <= \$11529_forever3163133\;
            when \$11529_forever3163133\ =>
              state_var7021 <= \$11529_forever3163133\;
            when \$11584_forever3163174\ =>
              state_var7021 <= \$11588_forever3163133\;
            when \$11588_forever3163133\ =>
              state_var7021 <= \$11588_forever3163133\;
            when \$11604_forever3163175\ =>
              state_var7021 <= \$11608_forever3163133\;
            when \$11608_forever3163133\ =>
              state_var7021 <= \$11608_forever3163133\;
            when \$11619_forever3163176\ =>
              state_var7021 <= \$11623_forever3163133\;
            when \$11623_forever3163133\ =>
              state_var7021 <= \$11623_forever3163133\;
            when \$11633_forever3163177\ =>
              state_var7021 <= \$11637_forever3163133\;
            when \$11637_forever3163133\ =>
              state_var7021 <= \$11637_forever3163133\;
            when \$11647_forever3163178\ =>
              state_var7021 <= \$11651_forever3163133\;
            when \$11651_forever3163133\ =>
              state_var7021 <= \$11651_forever3163133\;
            when \$11683_forever3163179\ =>
              state_var7021 <= \$11687_forever3163133\;
            when \$11687_forever3163133\ =>
              state_var7021 <= \$11687_forever3163133\;
            when \$11698_forever3163180\ =>
              state_var7021 <= \$11702_forever3163133\;
            when \$11702_forever3163133\ =>
              state_var7021 <= \$11702_forever3163133\;
            when \$11720_forever3163181\ =>
              state_var7021 <= \$11724_forever3163133\;
            when \$11724_forever3163133\ =>
              state_var7021 <= \$11724_forever3163133\;
            when \$11764_forever3163182\ =>
              state_var7021 <= \$11768_forever3163133\;
            when \$11768_forever3163133\ =>
              state_var7021 <= \$11768_forever3163133\;
            when \$11779_forever3163183\ =>
              state_var7021 <= \$11783_forever3163133\;
            when \$11783_forever3163133\ =>
              state_var7021 <= \$11783_forever3163133\;
            when \$11793_forever3163184\ =>
              state_var7021 <= \$11797_forever3163133\;
            when \$11797_forever3163133\ =>
              state_var7021 <= \$11797_forever3163133\;
            when \$11834_forever3163185\ =>
              state_var7021 <= \$11838_forever3163133\;
            when \$11838_forever3163133\ =>
              state_var7021 <= \$11838_forever3163133\;
            when \$11867_forever3163186\ =>
              state_var7021 <= \$11871_forever3163133\;
            when \$11871_forever3163133\ =>
              state_var7021 <= \$11871_forever3163133\;
            when \$11881_forever3163187\ =>
              state_var7021 <= \$11885_forever3163133\;
            when \$11885_forever3163133\ =>
              state_var7021 <= \$11885_forever3163133\;
            when \$11895_forever3163188\ =>
              state_var7021 <= \$11899_forever3163133\;
            when \$11899_forever3163133\ =>
              state_var7021 <= \$11899_forever3163133\;
            when \$11933_forever3163189\ =>
              state_var7021 <= \$11937_forever3163133\;
            when \$11937_forever3163133\ =>
              state_var7021 <= \$11937_forever3163133\;
            when \$11951_forever3163190\ =>
              state_var7021 <= \$11955_forever3163133\;
            when \$11955_forever3163133\ =>
              state_var7021 <= \$11955_forever3163133\;
            when \$11992_forever3163191\ =>
              state_var7021 <= \$11996_forever3163133\;
            when \$11996_forever3163133\ =>
              state_var7021 <= \$11996_forever3163133\;
            when \$12006_forever3163192\ =>
              state_var7021 <= \$12010_forever3163133\;
            when \$12010_forever3163133\ =>
              state_var7021 <= \$12010_forever3163133\;
            when \$12020_forever3163193\ =>
              state_var7021 <= \$12024_forever3163133\;
            when \$12024_forever3163133\ =>
              state_var7021 <= \$12024_forever3163133\;
            when \$12061_forever3163194\ =>
              state_var7021 <= \$12065_forever3163133\;
            when \$12065_forever3163133\ =>
              state_var7021 <= \$12065_forever3163133\;
            when \$12075_forever3163195\ =>
              state_var7021 <= \$12079_forever3163133\;
            when \$12079_forever3163133\ =>
              state_var7021 <= \$12079_forever3163133\;
            when \$12089_forever3163196\ =>
              state_var7021 <= \$12093_forever3163133\;
            when \$12093_forever3163133\ =>
              state_var7021 <= \$12093_forever3163133\;
            when \$12130_forever3163197\ =>
              state_var7021 <= \$12134_forever3163133\;
            when \$12134_forever3163133\ =>
              state_var7021 <= \$12134_forever3163133\;
            when \$12144_forever3163198\ =>
              state_var7021 <= \$12148_forever3163133\;
            when \$12148_forever3163133\ =>
              state_var7021 <= \$12148_forever3163133\;
            when \$12158_forever3163199\ =>
              state_var7021 <= \$12162_forever3163133\;
            when \$12162_forever3163133\ =>
              state_var7021 <= \$12162_forever3163133\;
            when \$12203_forever3163200\ =>
              state_var7021 <= \$12207_forever3163133\;
            when \$12207_forever3163133\ =>
              state_var7021 <= \$12207_forever3163133\;
            when \$12217_forever3163201\ =>
              state_var7021 <= \$12221_forever3163133\;
            when \$12221_forever3163133\ =>
              state_var7021 <= \$12221_forever3163133\;
            when \$12240_forever3163202\ =>
              state_var7021 <= \$12244_forever3163133\;
            when \$12244_forever3163133\ =>
              state_var7021 <= \$12244_forever3163133\;
            when \$12253_forever3163203\ =>
              state_var7021 <= \$12257_forever3163133\;
            when \$12257_forever3163133\ =>
              state_var7021 <= \$12257_forever3163133\;
            when \$12267_forever3163204\ =>
              state_var7021 <= \$12271_forever3163133\;
            when \$12271_forever3163133\ =>
              state_var7021 <= \$12271_forever3163133\;
            when \$12281_forever3163205\ =>
              state_var7021 <= \$12285_forever3163133\;
            when \$12285_forever3163133\ =>
              state_var7021 <= \$12285_forever3163133\;
            when \$12326_forever3163206\ =>
              state_var7021 <= \$12330_forever3163133\;
            when \$12330_forever3163133\ =>
              state_var7021 <= \$12330_forever3163133\;
            when \$12340_forever3163207\ =>
              state_var7021 <= \$12344_forever3163133\;
            when \$12344_forever3163133\ =>
              state_var7021 <= \$12344_forever3163133\;
            when \$12363_forever3163208\ =>
              state_var7021 <= \$12367_forever3163133\;
            when \$12367_forever3163133\ =>
              state_var7021 <= \$12367_forever3163133\;
            when \$12376_forever3163209\ =>
              state_var7021 <= \$12380_forever3163133\;
            when \$12380_forever3163133\ =>
              state_var7021 <= \$12380_forever3163133\;
            when \$12390_forever3163210\ =>
              state_var7021 <= \$12394_forever3163133\;
            when \$12394_forever3163133\ =>
              state_var7021 <= \$12394_forever3163133\;
            when \$12404_forever3163211\ =>
              state_var7021 <= \$12408_forever3163133\;
            when \$12408_forever3163133\ =>
              state_var7021 <= \$12408_forever3163133\;
            when \$12449_forever3163212\ =>
              state_var7021 <= \$12453_forever3163133\;
            when \$12453_forever3163133\ =>
              state_var7021 <= \$12453_forever3163133\;
            when \$12463_forever3163213\ =>
              state_var7021 <= \$12467_forever3163133\;
            when \$12467_forever3163133\ =>
              state_var7021 <= \$12467_forever3163133\;
            when \$12486_forever3163214\ =>
              state_var7021 <= \$12490_forever3163133\;
            when \$12490_forever3163133\ =>
              state_var7021 <= \$12490_forever3163133\;
            when \$12499_forever3163215\ =>
              state_var7021 <= \$12503_forever3163133\;
            when \$12503_forever3163133\ =>
              state_var7021 <= \$12503_forever3163133\;
            when \$12513_forever3163216\ =>
              state_var7021 <= \$12517_forever3163133\;
            when \$12517_forever3163133\ =>
              state_var7021 <= \$12517_forever3163133\;
            when \$12527_forever3163217\ =>
              state_var7021 <= \$12531_forever3163133\;
            when \$12531_forever3163133\ =>
              state_var7021 <= \$12531_forever3163133\;
            when \$12573_forever3163218\ =>
              state_var7021 <= \$12577_forever3163133\;
            when \$12577_forever3163133\ =>
              state_var7021 <= \$12577_forever3163133\;
            when \$12621_forever3163219\ =>
              state_var7021 <= \$12625_forever3163133\;
            when \$12625_forever3163133\ =>
              state_var7021 <= \$12625_forever3163133\;
            when \$12634_forever3163220\ =>
              state_var7021 <= \$12638_forever3163133\;
            when \$12638_forever3163133\ =>
              state_var7021 <= \$12638_forever3163133\;
            when \$12648_forever3163221\ =>
              state_var7021 <= \$12652_forever3163133\;
            when \$12652_forever3163133\ =>
              state_var7021 <= \$12652_forever3163133\;
            when \$12662_forever3163222\ =>
              state_var7021 <= \$12666_forever3163133\;
            when \$12666_forever3163133\ =>
              state_var7021 <= \$12666_forever3163133\;
            when \$12707_forever3163223\ =>
              state_var7021 <= \$12711_forever3163133\;
            when \$12711_forever3163133\ =>
              state_var7021 <= \$12711_forever3163133\;
            when \$12723_forever3163225\ =>
              state_var7021 <= \$12727_forever3163133\;
            when \$12727_forever3163133\ =>
              state_var7021 <= \$12727_forever3163133\;
            when \$12734_forever3163224\ =>
              state_var7021 <= \$12738_forever3163133\;
            when \$12738_forever3163133\ =>
              state_var7021 <= \$12738_forever3163133\;
            when \$12747_forever3163226\ =>
              state_var7021 <= \$12751_forever3163133\;
            when \$12751_forever3163133\ =>
              state_var7021 <= \$12751_forever3163133\;
            when \$12761_forever3163227\ =>
              state_var7021 <= \$12765_forever3163133\;
            when \$12765_forever3163133\ =>
              state_var7021 <= \$12765_forever3163133\;
            when \$12806_forever3163228\ =>
              state_var7021 <= \$12810_forever3163133\;
            when \$12810_forever3163133\ =>
              state_var7021 <= \$12810_forever3163133\;
            when \$12820_forever3163229\ =>
              state_var7021 <= \$12824_forever3163133\;
            when \$12824_forever3163133\ =>
              state_var7021 <= \$12824_forever3163133\;
            when \$12834_forever3163230\ =>
              state_var7021 <= \$12838_forever3163133\;
            when \$12838_forever3163133\ =>
              state_var7021 <= \$12838_forever3163133\;
            when \$12847_forever3163231\ =>
              state_var7021 <= \$12851_forever3163133\;
            when \$12851_forever3163133\ =>
              state_var7021 <= \$12851_forever3163133\;
            when \$12861_forever3163232\ =>
              state_var7021 <= \$12865_forever3163133\;
            when \$12865_forever3163133\ =>
              state_var7021 <= \$12865_forever3163133\;
            when \$12906_forever3163233\ =>
              state_var7021 <= \$12910_forever3163133\;
            when \$12910_forever3163133\ =>
              state_var7021 <= \$12910_forever3163133\;
            when \$12920_forever3163234\ =>
              state_var7021 <= \$12924_forever3163133\;
            when \$12924_forever3163133\ =>
              state_var7021 <= \$12924_forever3163133\;
            when \$12934_forever3163235\ =>
              state_var7021 <= \$12938_forever3163133\;
            when \$12938_forever3163133\ =>
              state_var7021 <= \$12938_forever3163133\;
            when \$12947_forever3163236\ =>
              state_var7021 <= \$12951_forever3163133\;
            when \$12951_forever3163133\ =>
              state_var7021 <= \$12951_forever3163133\;
            when \$12961_forever3163237\ =>
              state_var7021 <= \$12965_forever3163133\;
            when \$12965_forever3163133\ =>
              state_var7021 <= \$12965_forever3163133\;
            when \$13006_forever3163238\ =>
              state_var7021 <= \$13010_forever3163133\;
            when \$13010_forever3163133\ =>
              state_var7021 <= \$13010_forever3163133\;
            when \$13020_forever3163239\ =>
              state_var7021 <= \$13024_forever3163133\;
            when \$13024_forever3163133\ =>
              state_var7021 <= \$13024_forever3163133\;
            when \$13034_forever3163240\ =>
              state_var7021 <= \$13038_forever3163133\;
            when \$13038_forever3163133\ =>
              state_var7021 <= \$13038_forever3163133\;
            when \$13047_forever3163241\ =>
              state_var7021 <= \$13051_forever3163133\;
            when \$13051_forever3163133\ =>
              state_var7021 <= \$13051_forever3163133\;
            when \$13061_forever3163242\ =>
              state_var7021 <= \$13065_forever3163133\;
            when \$13065_forever3163133\ =>
              state_var7021 <= \$13065_forever3163133\;
            when \$13106_forever3163243\ =>
              state_var7021 <= \$13110_forever3163133\;
            when \$13110_forever3163133\ =>
              state_var7021 <= \$13110_forever3163133\;
            when \$13120_forever3163244\ =>
              state_var7021 <= \$13124_forever3163133\;
            when \$13124_forever3163133\ =>
              state_var7021 <= \$13124_forever3163133\;
            when \$13134_forever3163245\ =>
              state_var7021 <= \$13138_forever3163133\;
            when \$13138_forever3163133\ =>
              state_var7021 <= \$13138_forever3163133\;
            when \$13147_forever3163246\ =>
              state_var7021 <= \$13151_forever3163133\;
            when \$13151_forever3163133\ =>
              state_var7021 <= \$13151_forever3163133\;
            when \$13161_forever3163247\ =>
              state_var7021 <= \$13165_forever3163133\;
            when \$13165_forever3163133\ =>
              state_var7021 <= \$13165_forever3163133\;
            when \$13194_forever3163248\ =>
              state_var7021 <= \$13198_forever3163133\;
            when \$13198_forever3163133\ =>
              state_var7021 <= \$13198_forever3163133\;
            when \$13206_forever3163249\ =>
              state_var7021 <= \$13210_forever3163133\;
            when \$13210_forever3163133\ =>
              state_var7021 <= \$13210_forever3163133\;
            when \$13242_forever3163250\ =>
              state_var7021 <= \$13246_forever3163133\;
            when \$13246_forever3163133\ =>
              state_var7021 <= \$13246_forever3163133\;
            when \$13257_forever3163251\ =>
              state_var7021 <= \$13261_forever3163133\;
            when \$13261_forever3163133\ =>
              state_var7021 <= \$13261_forever3163133\;
            when \$13270_forever3163252\ =>
              state_var7021 <= \$13274_forever3163133\;
            when \$13274_forever3163133\ =>
              state_var7021 <= \$13274_forever3163133\;
            when \$13283_forever3163253\ =>
              state_var7021 <= \$13287_forever3163133\;
            when \$13287_forever3163133\ =>
              state_var7021 <= \$13287_forever3163133\;
            when \$13305_forever3163254\ =>
              state_var7021 <= \$13309_forever3163133\;
            when \$13309_forever3163133\ =>
              state_var7021 <= \$13309_forever3163133\;
            when \$13318_list_tail2653256\ =>
              \$v5284\ := eclat_lt(X"0000000" & X"0" & \$13318_list_tail2653256_arg\(36 to 67));
              if \$v5284\(0) = '1' then
                \$v5282\ := \$13318_list_tail2653256_arg\(0 to 35);
                \$v5283\ := \$v5282\(0 to 3);
                \$v5277\ := \$v5282\(4 to 35);
                case \$v5283\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13339_forever3163255\;
                when "0000" =>
                  \$13347_i\ := \$v5277\(0 to 31);
                  \$v5281\ := \$$10696_ram_ptr_take\;
                  if \$v5281\(0) = '1' then
                    state_var7021 <= q_wait5280;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$13347_i\));
                    state_var7021 <= pause_getI5278;
                  end if;
                when others =>
                  
                end case;
              else
                \$13318_list_tail2653256_result\ := \$13318_list_tail2653256_arg\(0 to 35);
                \$13295\ := \$13318_list_tail2653256_result\;
                \$v5275\ := \$13295\;
                \$v5276\ := \$v5275\(0 to 3);
                \$v5270\ := \$v5275\(4 to 35);
                case \$v5276\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13305_forever3163254\;
                when "0000" =>
                  \$13313_i\ := \$v5270\(0 to 31);
                  \$v5274\ := \$$10696_ram_ptr_take\;
                  if \$v5274\(0) = '1' then
                    state_var7021 <= q_wait5273;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$13313_i\));
                    state_var7021 <= pause_getI5271;
                  end if;
                when others =>
                  
                end case;
              end if;
            when \$13339_forever3163255\ =>
              state_var7021 <= \$13343_forever3163133\;
            when \$13343_forever3163133\ =>
              state_var7021 <= \$13343_forever3163133\;
            when \$13360_forever3163257\ =>
              state_var7021 <= \$13364_forever3163133\;
            when \$13364_forever3163133\ =>
              state_var7021 <= \$13364_forever3163133\;
            when \$13374_forever3163258\ =>
              state_var7021 <= \$13378_forever3163133\;
            when \$13378_forever3163133\ =>
              state_var7021 <= \$13378_forever3163133\;
            when \$13388_forever3163259\ =>
              state_var7021 <= \$13392_forever3163133\;
            when \$13392_forever3163133\ =>
              state_var7021 <= \$13392_forever3163133\;
            when \$13420_forever3163260\ =>
              state_var7021 <= \$13424_forever3163133\;
            when \$13424_forever3163133\ =>
              state_var7021 <= \$13424_forever3163133\;
            when \$13434_forever3163261\ =>
              state_var7021 <= \$13438_forever3163133\;
            when \$13438_forever3163133\ =>
              state_var7021 <= \$13438_forever3163133\;
            when \$13451_forever3163262\ =>
              state_var7021 <= \$13455_forever3163133\;
            when \$13455_forever3163133\ =>
              state_var7021 <= \$13455_forever3163133\;
            when \$13474_forever3163263\ =>
              state_var7021 <= \$13478_forever3163133\;
            when \$13478_forever3163133\ =>
              state_var7021 <= \$13478_forever3163133\;
            when \$13487_forever3163264\ =>
              state_var7021 <= \$13491_forever3163133\;
            when \$13491_forever3163133\ =>
              state_var7021 <= \$13491_forever3163133\;
            when \$13500_list_tail2653266\ =>
              \$v5365\ := eclat_lt(X"0000000" & X"0" & \$13500_list_tail2653266_arg\(36 to 67));
              if \$v5365\(0) = '1' then
                \$v5363\ := \$13500_list_tail2653266_arg\(0 to 35);
                \$v5364\ := \$v5363\(0 to 3);
                \$v5358\ := \$v5363\(4 to 35);
                case \$v5364\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13521_forever3163265\;
                when "0000" =>
                  \$13529_i\ := \$v5358\(0 to 31);
                  \$v5362\ := \$$10696_ram_ptr_take\;
                  if \$v5362\(0) = '1' then
                    state_var7021 <= q_wait5361;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$13529_i\));
                    state_var7021 <= pause_getI5359;
                  end if;
                when others =>
                  
                end case;
              else
                \$13500_list_tail2653266_result\ := \$13500_list_tail2653266_arg\(0 to 35);
                \$13446\ := \$13500_list_tail2653266_result\;
                \$v5356\ := \$13446\;
                \$v5357\ := \$v5356\(0 to 3);
                \$v5337\ := \$v5356\(4 to 35);
                case \$v5357\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't field0_set"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13451_forever3163262\;
                when "0000" =>
                  \$13459_i\ := \$v5337\(0 to 31);
                  \$v5354\ := \$13446\;
                  \$v5355\ := \$v5354\(0 to 3);
                  \$v5349\ := \$v5354\(4 to 35);
                  case \$v5355\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$13487_forever3163264\;
                  when "0000" =>
                    \$13495_i\ := \$v5349\(0 to 31);
                    \$v5353\ := \$$10696_ram_ptr_take\;
                    if \$v5353\(0) = '1' then
                      state_var7021 <= q_wait5352;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$13495_i\));
                      state_var7021 <= pause_getI5350;
                    end if;
                  when others =>
                    
                  end case;
                when others =>
                  
                end case;
              end if;
            when \$13521_forever3163265\ =>
              state_var7021 <= \$13525_forever3163133\;
            when \$13525_forever3163133\ =>
              state_var7021 <= \$13525_forever3163133\;
            when \$13537_forever3163267\ =>
              state_var7021 <= \$13541_forever3163133\;
            when \$13541_forever3163133\ =>
              state_var7021 <= \$13541_forever3163133\;
            when \$13560_forever3163268\ =>
              state_var7021 <= \$13564_forever3163133\;
            when \$13564_forever3163133\ =>
              state_var7021 <= \$13564_forever3163133\;
            when \$13573_forever3163269\ =>
              state_var7021 <= \$13577_forever3163133\;
            when \$13577_forever3163133\ =>
              state_var7021 <= \$13577_forever3163133\;
            when \$13587_forever3163270\ =>
              state_var7021 <= \$13591_forever3163133\;
            when \$13591_forever3163133\ =>
              state_var7021 <= \$13591_forever3163133\;
            when \$13618_forever3163271\ =>
              state_var7021 <= \$13622_forever3163133\;
            when \$13622_forever3163133\ =>
              state_var7021 <= \$13622_forever3163133\;
            when \$13632_forever3163272\ =>
              state_var7021 <= \$13636_forever3163133\;
            when \$13636_forever3163133\ =>
              state_var7021 <= \$13636_forever3163133\;
            when \$13653_forever3163273\ =>
              state_var7021 <= \$13657_forever3163133\;
            when \$13657_forever3163133\ =>
              state_var7021 <= \$13657_forever3163133\;
            when \$13676_forever3163274\ =>
              state_var7021 <= \$13680_forever3163133\;
            when \$13680_forever3163133\ =>
              state_var7021 <= \$13680_forever3163133\;
            when \$13689_list_tail2653276\ =>
              \$v5483\ := eclat_lt(X"0000000" & X"0" & \$13689_list_tail2653276_arg\(36 to 67));
              if \$v5483\(0) = '1' then
                \$v5481\ := \$13689_list_tail2653276_arg\(0 to 35);
                \$v5482\ := \$v5481\(0 to 3);
                \$v5476\ := \$v5481\(4 to 35);
                case \$v5482\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13710_forever3163275\;
                when "0000" =>
                  \$13718_i\ := \$v5476\(0 to 31);
                  \$v5480\ := \$$10696_ram_ptr_take\;
                  if \$v5480\(0) = '1' then
                    state_var7021 <= q_wait5479;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$13718_i\));
                    state_var7021 <= pause_getI5477;
                  end if;
                when others =>
                  
                end case;
              else
                \$13689_list_tail2653276_result\ := \$13689_list_tail2653276_arg\(0 to 35);
                \$13666\ := \$13689_list_tail2653276_result\;
                \$v5474\ := \$13666\;
                \$v5475\ := \$v5474\(0 to 3);
                \$v5469\ := \$v5474\(4 to 35);
                case \$v5475\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13676_forever3163274\;
                when "0000" =>
                  \$13684_i\ := \$v5469\(0 to 31);
                  \$v5473\ := \$$10696_ram_ptr_take\;
                  if \$v5473\(0) = '1' then
                    state_var7021 <= q_wait5472;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$13684_i\));
                    state_var7021 <= pause_getI5470;
                  end if;
                when others =>
                  
                end case;
              end if;
            when \$13710_forever3163275\ =>
              state_var7021 <= \$13714_forever3163133\;
            when \$13714_forever3163133\ =>
              state_var7021 <= \$13714_forever3163133\;
            when \$13731_forever3163277\ =>
              state_var7021 <= \$13735_forever3163133\;
            when \$13735_forever3163133\ =>
              state_var7021 <= \$13735_forever3163133\;
            when \$13761_forever3163278\ =>
              state_var7021 <= \$13765_forever3163133\;
            when \$13765_forever3163133\ =>
              state_var7021 <= \$13765_forever3163133\;
            when \$13775_forever3163279\ =>
              state_var7021 <= \$13779_forever3163133\;
            when \$13779_forever3163133\ =>
              state_var7021 <= \$13779_forever3163133\;
            when \$13796_forever3163280\ =>
              state_var7021 <= \$13800_forever3163133\;
            when \$13800_forever3163133\ =>
              state_var7021 <= \$13800_forever3163133\;
            when \$13821_forever3163281\ =>
              state_var7021 <= \$13825_forever3163133\;
            when \$13825_forever3163133\ =>
              state_var7021 <= \$13825_forever3163133\;
            when \$13842_forever3163282\ =>
              state_var7021 <= \$13846_forever3163133\;
            when \$13846_forever3163133\ =>
              state_var7021 <= \$13846_forever3163133\;
            when \$13856_forever3163283\ =>
              state_var7021 <= \$13860_forever3163133\;
            when \$13860_forever3163133\ =>
              state_var7021 <= \$13860_forever3163133\;
            when \$13878_forever3163284\ =>
              state_var7021 <= \$13882_forever3163133\;
            when \$13882_forever3163133\ =>
              state_var7021 <= \$13882_forever3163133\;
            when \$13892_forever3163134\ =>
              state_var7021 <= \$13896_forever3163133\;
            when \$13896_forever3163133\ =>
              state_var7021 <= \$13896_forever3163133\;
            when \$13905_forever3163285\ =>
              state_var7021 <= \$13909_forever3163133\;
            when \$13909_forever3163133\ =>
              state_var7021 <= \$13909_forever3163133\;
            when \$13931_forever3163286\ =>
              state_var7021 <= \$13935_forever3163133\;
            when \$13935_forever3163133\ =>
              state_var7021 <= \$13935_forever3163133\;
            when \$13950_forever3163287\ =>
              state_var7021 <= \$13954_forever3163133\;
            when \$13954_forever3163133\ =>
              state_var7021 <= \$13954_forever3163133\;
            when \$13977_forever3163288\ =>
              state_var7021 <= \$13981_forever3163133\;
            when \$13981_forever3163133\ =>
              state_var7021 <= \$13981_forever3163133\;
            when \$13991_forever3163289\ =>
              state_var7021 <= \$13995_forever3163133\;
            when \$13995_forever3163133\ =>
              state_var7021 <= \$13995_forever3163133\;
            when \$14004_forever3163290\ =>
              state_var7021 <= \$14008_forever3163133\;
            when \$14008_forever3163133\ =>
              state_var7021 <= \$14008_forever3163133\;
            when \$14037_forever3163291\ =>
              state_var7021 <= \$14041_forever3163133\;
            when \$14041_forever3163133\ =>
              state_var7021 <= \$14041_forever3163133\;
            when \$14050_forever3163292\ =>
              state_var7021 <= \$14054_forever3163133\;
            when \$14054_forever3163133\ =>
              state_var7021 <= \$14054_forever3163133\;
            when \$14064_forever3163293\ =>
              state_var7021 <= \$14068_forever3163133\;
            when \$14068_forever3163133\ =>
              state_var7021 <= \$14068_forever3163133\;
            when \$14090_forever3163294\ =>
              state_var7021 <= \$14094_forever3163133\;
            when \$14094_forever3163133\ =>
              state_var7021 <= \$14094_forever3163133\;
            when \$14104_forever3163295\ =>
              state_var7021 <= \$14108_forever3163133\;
            when \$14108_forever3163133\ =>
              state_var7021 <= \$14108_forever3163133\;
            when \$14117_forever3163296\ =>
              state_var7021 <= \$14121_forever3163133\;
            when \$14121_forever3163133\ =>
              state_var7021 <= \$14121_forever3163133\;
            when \$14150_forever3163297\ =>
              state_var7021 <= \$14154_forever3163133\;
            when \$14154_forever3163133\ =>
              state_var7021 <= \$14154_forever3163133\;
            when \$14163_forever3163298\ =>
              state_var7021 <= \$14167_forever3163133\;
            when \$14167_forever3163133\ =>
              state_var7021 <= \$14167_forever3163133\;
            when \$14177_forever3163299\ =>
              state_var7021 <= \$14181_forever3163133\;
            when \$14181_forever3163133\ =>
              state_var7021 <= \$14181_forever3163133\;
            when \$14203_forever3163300\ =>
              state_var7021 <= \$14207_forever3163133\;
            when \$14207_forever3163133\ =>
              state_var7021 <= \$14207_forever3163133\;
            when \$14217_forever3163301\ =>
              state_var7021 <= \$14221_forever3163133\;
            when \$14221_forever3163133\ =>
              state_var7021 <= \$14221_forever3163133\;
            when \$14230_forever3163302\ =>
              state_var7021 <= \$14234_forever3163133\;
            when \$14234_forever3163133\ =>
              state_var7021 <= \$14234_forever3163133\;
            when \$14263_forever3163303\ =>
              state_var7021 <= \$14267_forever3163133\;
            when \$14267_forever3163133\ =>
              state_var7021 <= \$14267_forever3163133\;
            when \$14276_forever3163304\ =>
              state_var7021 <= \$14280_forever3163133\;
            when \$14280_forever3163133\ =>
              state_var7021 <= \$14280_forever3163133\;
            when \$14290_forever3163305\ =>
              state_var7021 <= \$14294_forever3163133\;
            when \$14294_forever3163133\ =>
              state_var7021 <= \$14294_forever3163133\;
            when \$14311_forever3163306\ =>
              state_var7021 <= \$14315_forever3163133\;
            when \$14315_forever3163133\ =>
              state_var7021 <= \$14315_forever3163133\;
            when \$14325_forever3163307\ =>
              state_var7021 <= \$14329_forever3163133\;
            when \$14329_forever3163133\ =>
              state_var7021 <= \$14329_forever3163133\;
            when \$14338_forever3163308\ =>
              state_var7021 <= \$14342_forever3163133\;
            when \$14342_forever3163133\ =>
              state_var7021 <= \$14342_forever3163133\;
            when \$14369_forever3163309\ =>
              state_var7021 <= \$14373_forever3163133\;
            when \$14373_forever3163133\ =>
              state_var7021 <= \$14373_forever3163133\;
            when \$14382_forever3163310\ =>
              state_var7021 <= \$14386_forever3163133\;
            when \$14386_forever3163133\ =>
              state_var7021 <= \$14386_forever3163133\;
            when \$14396_forever3163311\ =>
              state_var7021 <= \$14400_forever3163133\;
            when \$14400_forever3163133\ =>
              state_var7021 <= \$14400_forever3163133\;
            when \$14423_forever3163312\ =>
              state_var7021 <= \$14427_forever3163133\;
            when \$14427_forever3163133\ =>
              state_var7021 <= \$14427_forever3163133\;
            when \$14437_forever3163313\ =>
              state_var7021 <= \$14441_forever3163133\;
            when \$14441_forever3163133\ =>
              state_var7021 <= \$14441_forever3163133\;
            when \$14450_forever3163314\ =>
              state_var7021 <= \$14454_forever3163133\;
            when \$14454_forever3163133\ =>
              state_var7021 <= \$14454_forever3163133\;
            when \$14464_forever3163315\ =>
              state_var7021 <= \$14468_forever3163133\;
            when \$14468_forever3163133\ =>
              state_var7021 <= \$14468_forever3163133\;
            when \$14481_decode_loop310\ =>
              \$v6436\ := \$$10701_pos_ptr_take\;
              if \$v6436\(0) = '1' then
                state_var7021 <= q_wait6435;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6433;
              end if;
            when \$14511_loop311\ =>
              \$v6424\ := eclat_lt(eclat_add(eclat_vector_get(X"000000" & X"14" & X"000000" & X"1e" & X"0000000" & X"0" & X"0000000" & X"a" & X"0000000" & X"b" & X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31),32) & X"0000000" & X"2") & \$14511_loop311_arg\(32 to 63));
              if \$v6424\(0) = '1' then
                \$14511_loop311_arg\ := eclat_add(\$14511_loop311_arg\(0 to 31) & X"0000000" & X"1") & eclat_sub(\$14511_loop311_arg\(32 to 63) & eclat_add(eclat_vector_get(X"000000" & X"14" & X"000000" & X"1e" & X"0000000" & X"0" & X"0000000" & X"a" & X"0000000" & X"b" & X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31),32) & X"0000000" & X"3")) & \$14511_loop311_arg\(64 to 95) & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
                state_var7021 <= \$14511_loop311\;
              else
                \$v6423\ := eclat_lt(X"000000" & X"5a" & \$14511_loop311_arg\(64 to 95));
                if \$v6423\(0) = '1' then
                  \$v6053\ := \$$10697_stack_ptr_take\;
                  if \$v6053\(0) = '1' then
                    state_var7021 <= q_wait6052;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI6050;
                  end if;
                else
                  \$v6422\ := eclat_eq(\$14511_loop311_arg\(0 to 31) & X"0000000" & X"0");
                  if \$v6422\(0) = '1' then
                    \$v6421\ := \$$10702_brk_ptr_take\;
                    if \$v6421\(0) = '1' then
                      state_var7021 <= q_wait6420;
                    else
                      \$$10702_brk_ptr_take\(0) := '1';
                      \$$10702_brk_ptr\ <= 0;
                      state_var7021 <= pause_getI6418;
                    end if;
                  else
                    \$v6378\ := eclat_lt(\$14511_loop311_arg\(32 to 63) & eclat_vector_get(X"000000" & X"14" & X"000000" & X"1e" & X"0000000" & X"0" & X"0000000" & X"a" & X"0000000" & X"b" & X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31),32));
                    if \$v6378\(0) = '1' then
                      \$v6331\ := eclat_lt(\$14511_loop311_arg\(0 to 31) & X"0000000" & X"3");
                      if \$v6331\(0) = '1' then
                        \$v6329\ := \$$10699_symtbl_ptr_take\;
                        if \$v6329\(0) = '1' then
                          state_var7021 <= q_wait6328;
                        else
                          \$$10699_symtbl_ptr_take\(0) := '1';
                          \$$10699_symtbl_ptr\ <= 0;
                          state_var7021 <= pause_getI6326;
                        end if;
                      else
                        \$v6330\ := \$14511_loop311_arg\(32 to 63);
                        \$14533_opnd\ := "0001" & \$v6330\;
                        \$v6310\ := eclat_lt(X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31));
                        if \$v6310\(0) = '1' then
                          \$v6235\ := \$$10697_stack_ptr_take\;
                          if \$v6235\(0) = '1' then
                            state_var7021 <= q_wait6234;
                          else
                            \$$10697_stack_ptr_take\(0) := '1';
                            \$$10697_stack_ptr\ <= 0;
                            state_var7021 <= pause_getI6232;
                          end if;
                        else
                          \$v6309\ := \$$10697_stack_ptr_take\;
                          if \$v6309\(0) = '1' then
                            state_var7021 <= q_wait6308;
                          else
                            \$$10697_stack_ptr_take\(0) := '1';
                            \$$10697_stack_ptr\ <= 0;
                            state_var7021 <= pause_getI6306;
                          end if;
                        end if;
                      end if;
                    else
                      \$v6377\ := eclat_eq(\$14511_loop311_arg\(32 to 63) & eclat_vector_get(X"000000" & X"14" & X"000000" & X"1e" & X"0000000" & X"0" & X"0000000" & X"a" & X"0000000" & X"b" & X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31),32));
                      if \$v6377\(0) = '1' then
                        \$14939_get_int268_arg\ := X"0000000" & X"0" & eclat_unit;
                        state_var7021 <= \$14939_get_int268\;
                      else
                        \$14897_get_int268_arg\ := eclat_sub(eclat_sub(\$14511_loop311_arg\(32 to 63) & eclat_vector_get(X"000000" & X"14" & X"000000" & X"1e" & X"0000000" & X"0" & X"0000000" & X"a" & X"0000000" & X"b" & X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31),32)) & X"0000000" & X"1") & eclat_unit;
                        state_var7021 <= \$14897_get_int268\;
                      end if;
                    end if;
                  end if;
                end if;
              end if;
            when \$14548_forever3163316\ =>
              state_var7021 <= \$14552_forever3163133\;
            when \$14552_forever3163133\ =>
              state_var7021 <= \$14552_forever3163133\;
            when \$14572_forever3163317\ =>
              state_var7021 <= \$14576_forever3163133\;
            when \$14576_forever3163133\ =>
              state_var7021 <= \$14576_forever3163133\;
            when \$14586_forever3163318\ =>
              state_var7021 <= \$14590_forever3163133\;
            when \$14590_forever3163133\ =>
              state_var7021 <= \$14590_forever3163133\;
            when \$14617_forever3163319\ =>
              state_var7021 <= \$14621_forever3163133\;
            when \$14621_forever3163133\ =>
              state_var7021 <= \$14621_forever3163133\;
            when \$14632_forever3163320\ =>
              state_var7021 <= \$14636_forever3163133\;
            when \$14636_forever3163133\ =>
              state_var7021 <= \$14636_forever3163133\;
            when \$14673_forever3163321\ =>
              state_var7021 <= \$14677_forever3163133\;
            when \$14677_forever3163133\ =>
              state_var7021 <= \$14677_forever3163133\;
            when \$14697_forever3163322\ =>
              state_var7021 <= \$14701_forever3163133\;
            when \$14701_forever3163133\ =>
              state_var7021 <= \$14701_forever3163133\;
            when \$14711_forever3163323\ =>
              state_var7021 <= \$14715_forever3163133\;
            when \$14715_forever3163133\ =>
              state_var7021 <= \$14715_forever3163133\;
            when \$14740_forever3163324\ =>
              state_var7021 <= \$14744_forever3163133\;
            when \$14744_forever3163133\ =>
              state_var7021 <= \$14744_forever3163133\;
            when \$14755_forever3163325\ =>
              state_var7021 <= \$14759_forever3163133\;
            when \$14759_forever3163133\ =>
              state_var7021 <= \$14759_forever3163133\;
            when \$14785_forever3163326\ =>
              state_var7021 <= \$14789_forever3163133\;
            when \$14789_forever3163133\ =>
              state_var7021 <= \$14789_forever3163133\;
            when \$14811_forever3163327\ =>
              state_var7021 <= \$14815_forever3163133\;
            when \$14815_forever3163133\ =>
              state_var7021 <= \$14815_forever3163133\;
            when \$14826_forever3163328\ =>
              state_var7021 <= \$14830_forever3163133\;
            when \$14830_forever3163133\ =>
              state_var7021 <= \$14830_forever3163133\;
            when \$14850_forever3163329\ =>
              state_var7021 <= \$14854_forever3163133\;
            when \$14854_forever3163133\ =>
              state_var7021 <= \$14854_forever3163133\;
            when \$14863_list_tail2653331\ =>
              \$v6359\ := eclat_lt(X"0000000" & X"0" & \$14863_list_tail2653331_arg\(36 to 67));
              if \$v6359\(0) = '1' then
                \$v6357\ := \$14863_list_tail2653331_arg\(0 to 35);
                \$v6358\ := \$v6357\(0 to 3);
                \$v6352\ := \$v6357\(4 to 35);
                case \$v6358\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14884_forever3163330\;
                when "0000" =>
                  \$14892_i\ := \$v6352\(0 to 31);
                  \$v6356\ := \$$10696_ram_ptr_take\;
                  if \$v6356\(0) = '1' then
                    state_var7021 <= q_wait6355;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14892_i\));
                    state_var7021 <= pause_getI6353;
                  end if;
                when others =>
                  
                end case;
              else
                \$14863_list_tail2653331_result\ := \$14863_list_tail2653331_arg\(0 to 35);
                \$14840\ := \$14863_list_tail2653331_result\;
                \$v6350\ := \$14840\;
                \$v6351\ := \$v6350\(0 to 3);
                \$v6345\ := \$v6350\(4 to 35);
                case \$v6351\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14850_forever3163329\;
                when "0000" =>
                  \$14858_i\ := \$v6345\(0 to 31);
                  \$v6349\ := \$$10696_ram_ptr_take\;
                  if \$v6349\(0) = '1' then
                    state_var7021 <= q_wait6348;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14858_i\));
                    state_var7021 <= pause_getI6346;
                  end if;
                when others =>
                  
                end case;
              end if;
            when \$14884_forever3163330\ =>
              state_var7021 <= \$14888_forever3163133\;
            when \$14888_forever3163133\ =>
              state_var7021 <= \$14888_forever3163133\;
            when \$14897_get_int268\ =>
              \$v6376\ := \$$10701_pos_ptr_take\;
              if \$v6376\(0) = '1' then
                state_var7021 <= q_wait6375;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6373;
              end if;
            when \$14939_get_int268\ =>
              \$v6344\ := \$$10701_pos_ptr_take\;
              if \$v6344\(0) = '1' then
                state_var7021 <= q_wait6343;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6341;
              end if;
            when \$14983_forever3163332\ =>
              state_var7021 <= \$14987_forever3163133\;
            when \$14987_forever3163133\ =>
              state_var7021 <= \$14987_forever3163133\;
            when \$14996_list_tail2653334\ =>
              \$v6325\ := eclat_lt(X"0000000" & X"0" & \$14996_list_tail2653334_arg\(36 to 67));
              if \$v6325\(0) = '1' then
                \$v6323\ := \$14996_list_tail2653334_arg\(0 to 35);
                \$v6324\ := \$v6323\(0 to 3);
                \$v6318\ := \$v6323\(4 to 35);
                case \$v6324\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$15017_forever3163333\;
                when "0000" =>
                  \$15025_i\ := \$v6318\(0 to 31);
                  \$v6322\ := \$$10696_ram_ptr_take\;
                  if \$v6322\(0) = '1' then
                    state_var7021 <= q_wait6321;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$15025_i\));
                    state_var7021 <= pause_getI6319;
                  end if;
                when others =>
                  
                end case;
              else
                \$14996_list_tail2653334_result\ := \$14996_list_tail2653334_arg\(0 to 35);
                \$14973\ := \$14996_list_tail2653334_result\;
                \$v6316\ := \$14973\;
                \$v6317\ := \$v6316\(0 to 3);
                \$v6311\ := \$v6316\(4 to 35);
                case \$v6317\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14983_forever3163332\;
                when "0000" =>
                  \$14991_i\ := \$v6311\(0 to 31);
                  \$v6315\ := \$$10696_ram_ptr_take\;
                  if \$v6315\(0) = '1' then
                    state_var7021 <= q_wait6314;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14991_i\));
                    state_var7021 <= pause_getI6312;
                  end if;
                when others =>
                  
                end case;
              end if;
            when \$15017_forever3163333\ =>
              state_var7021 <= \$15021_forever3163133\;
            when \$15021_forever3163133\ =>
              state_var7021 <= \$15021_forever3163133\;
            when \$15051_forever3163335\ =>
              state_var7021 <= \$15055_forever3163133\;
            when \$15055_forever3163133\ =>
              state_var7021 <= \$15055_forever3163133\;
            when \$15082_forever3163336\ =>
              state_var7021 <= \$15086_forever3163133\;
            when \$15086_forever3163133\ =>
              state_var7021 <= \$15086_forever3163133\;
            when \$15106_forever3163337\ =>
              state_var7021 <= \$15110_forever3163133\;
            when \$15110_forever3163133\ =>
              state_var7021 <= \$15110_forever3163133\;
            when \$15120_forever3163338\ =>
              state_var7021 <= \$15124_forever3163133\;
            when \$15124_forever3163133\ =>
              state_var7021 <= \$15124_forever3163133\;
            when \$15149_forever3163339\ =>
              state_var7021 <= \$15153_forever3163133\;
            when \$15153_forever3163133\ =>
              state_var7021 <= \$15153_forever3163133\;
            when \$15164_forever3163340\ =>
              state_var7021 <= \$15168_forever3163133\;
            when \$15168_forever3163133\ =>
              state_var7021 <= \$15168_forever3163133\;
            when \$15178_forever3163341\ =>
              state_var7021 <= \$15182_forever3163133\;
            when \$15182_forever3163133\ =>
              state_var7021 <= \$15182_forever3163133\;
            when \$15217_loop1312\ =>
              \$v6981\ := eclat_lt(X"0000000" & X"0" & \$15217_loop1312_arg\(0 to 31));
              if \$v6981\(0) = '1' then
                \$v6599\ := \$$10699_symtbl_ptr_take\;
                if \$v6599\(0) = '1' then
                  state_var7021 <= q_wait6598;
                else
                  \$$10699_symtbl_ptr_take\(0) := '1';
                  \$$10699_symtbl_ptr\ <= 0;
                  state_var7021 <= pause_getI6596;
                end if;
              else
                \$v6980\ := X"0000000" & X"0";
                \$15240_loop23133355_arg\ := "0000" & \$v6980\ & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
                state_var7021 <= \$15240_loop23133355\;
              end if;
            when \$15240_loop23133355\ =>
              \$v6979\ := \$$10701_pos_ptr_take\;
              if \$v6979\(0) = '1' then
                state_var7021 <= q_wait6978;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6976;
              end if;
            when \$15282_forever3163342\ =>
              state_var7021 <= \$15286_forever3163133\;
            when \$15286_forever3163133\ =>
              state_var7021 <= \$15286_forever3163133\;
            when \$15332_forever3163343\ =>
              state_var7021 <= \$15336_forever3163133\;
            when \$15336_forever3163133\ =>
              state_var7021 <= \$15336_forever3163133\;
            when \$15355_forever3163344\ =>
              state_var7021 <= \$15359_forever3163133\;
            when \$15359_forever3163133\ =>
              state_var7021 <= \$15359_forever3163133\;
            when \$15378_forever3163345\ =>
              state_var7021 <= \$15382_forever3163133\;
            when \$15382_forever3163133\ =>
              state_var7021 <= \$15382_forever3163133\;
            when \$15391_len_aux3143348\ =>
              \$v6917\ := \$15391_len_aux3143348_arg\(0 to 35);
              \$v6918\ := \$v6917\(0 to 3);
              \$v6916\ := \$v6917\(4 to 35);
              case \$v6918\ is
              when "0001" =>
                \$15399\ := eclat_false;
              when "0000" =>
                \$15449_i\ := \$v6916\(0 to 31);
                \$15399\ := eclat_if(eclat_ge(\$15449_i\ & X"0000000" & X"0") & eclat_lt(\$15449_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v6915\ := \$15399\;
              if \$v6915\(0) = '1' then
                \$v6913\ := \$15391_len_aux3143348_arg\(0 to 35);
                \$v6914\ := \$v6913\(0 to 3);
                \$v6908\ := \$v6913\(4 to 35);
                case \$v6914\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$15439_forever3163347\;
                when "0000" =>
                  \$15447_i\ := \$v6908\(0 to 31);
                  \$v6912\ := \$$10696_ram_ptr_take\;
                  if \$v6912\(0) = '1' then
                    state_var7021 <= q_wait6911;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$15447_i\));
                    state_var7021 <= pause_getI6909;
                  end if;
                when others =>
                  
                end case;
              else
                \$15400\ := eclat_false;
                \$v6896\ := \$15400\;
                if \$v6896\(0) = '1' then
                  \$v6894\ := \$15391_len_aux3143348_arg\(0 to 35);
                  \$v6895\ := \$v6894\(0 to 3);
                  \$v6889\ := \$v6894\(4 to 35);
                  case \$v6895\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15413_forever3163346\;
                  when "0000" =>
                    \$15421_i\ := \$v6889\(0 to 31);
                    \$v6893\ := \$$10696_ram_ptr_take\;
                    if \$v6893\(0) = '1' then
                      state_var7021 <= q_wait6892;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15421_i\));
                      state_var7021 <= pause_getI6890;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15391_len_aux3143348_result\ := \$15391_len_aux3143348_arg\(36 to 67);
                  \$15294\ := \$15391_len_aux3143348_result\;
                  \$v6888\ := \$$10702_brk_ptr_take\;
                  if \$v6888\(0) = '1' then
                    state_var7021 <= q_wait6887;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6885;
                  end if;
                end if;
              end if;
            when \$15413_forever3163346\ =>
              state_var7021 <= \$15417_forever3163133\;
            when \$15417_forever3163133\ =>
              state_var7021 <= \$15417_forever3163133\;
            when \$15439_forever3163347\ =>
              state_var7021 <= \$15443_forever3163133\;
            when \$15443_forever3163133\ =>
              state_var7021 <= \$15443_forever3163133\;
            when \$15496_forever3163349\ =>
              state_var7021 <= \$15500_forever3163133\;
            when \$15500_forever3163133\ =>
              state_var7021 <= \$15500_forever3163133\;
            when \$15519_forever3163350\ =>
              state_var7021 <= \$15523_forever3163133\;
            when \$15523_forever3163133\ =>
              state_var7021 <= \$15523_forever3163133\;
            when \$15542_forever3163351\ =>
              state_var7021 <= \$15546_forever3163133\;
            when \$15546_forever3163133\ =>
              state_var7021 <= \$15546_forever3163133\;
            when \$15555_len_aux3143354\ =>
              \$v6756\ := \$15555_len_aux3143354_arg\(0 to 35);
              \$v6757\ := \$v6756\(0 to 3);
              \$v6755\ := \$v6756\(4 to 35);
              case \$v6757\ is
              when "0001" =>
                \$15563\ := eclat_false;
              when "0000" =>
                \$15613_i\ := \$v6755\(0 to 31);
                \$15563\ := eclat_if(eclat_ge(\$15613_i\ & X"0000000" & X"0") & eclat_lt(\$15613_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v6754\ := \$15563\;
              if \$v6754\(0) = '1' then
                \$v6752\ := \$15555_len_aux3143354_arg\(0 to 35);
                \$v6753\ := \$v6752\(0 to 3);
                \$v6747\ := \$v6752\(4 to 35);
                case \$v6753\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$15603_forever3163353\;
                when "0000" =>
                  \$15611_i\ := \$v6747\(0 to 31);
                  \$v6751\ := \$$10696_ram_ptr_take\;
                  if \$v6751\(0) = '1' then
                    state_var7021 <= q_wait6750;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$15611_i\));
                    state_var7021 <= pause_getI6748;
                  end if;
                when others =>
                  
                end case;
              else
                \$15564\ := eclat_false;
                \$v6735\ := \$15564\;
                if \$v6735\(0) = '1' then
                  \$v6733\ := \$15555_len_aux3143354_arg\(0 to 35);
                  \$v6734\ := \$v6733\(0 to 3);
                  \$v6728\ := \$v6733\(4 to 35);
                  case \$v6734\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15577_forever3163352\;
                  when "0000" =>
                    \$15585_i\ := \$v6728\(0 to 31);
                    \$v6732\ := \$$10696_ram_ptr_take\;
                    if \$v6732\(0) = '1' then
                      state_var7021 <= q_wait6731;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15585_i\));
                      state_var7021 <= pause_getI6729;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15555_len_aux3143354_result\ := \$15555_len_aux3143354_arg\(36 to 67);
                  \$15455\ := \$15555_len_aux3143354_result\;
                  \$v6727\ := \$$10702_brk_ptr_take\;
                  if \$v6727\(0) = '1' then
                    state_var7021 <= q_wait6726;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6724;
                  end if;
                end if;
              end if;
            when \$15577_forever3163352\ =>
              state_var7021 <= \$15581_forever3163133\;
            when \$15581_forever3163133\ =>
              state_var7021 <= \$15581_forever3163133\;
            when \$15603_forever3163353\ =>
              state_var7021 <= \$15607_forever3163133\;
            when \$15607_forever3163133\ =>
              state_var7021 <= \$15607_forever3163133\;
            when \$15663_forever3163356\ =>
              state_var7021 <= \$15667_forever3163133\;
            when \$15667_forever3163133\ =>
              state_var7021 <= \$15667_forever3163133\;
            when \$15686_forever3163357\ =>
              state_var7021 <= \$15690_forever3163133\;
            when \$15690_forever3163133\ =>
              state_var7021 <= \$15690_forever3163133\;
            when \$15710_forever3163358\ =>
              state_var7021 <= \$15714_forever3163133\;
            when \$15714_forever3163133\ =>
              state_var7021 <= \$15714_forever3163133\;
            when \$15724_len_aux3143361\ =>
              \$v6593\ := \$15724_len_aux3143361_arg\(0 to 35);
              \$v6594\ := \$v6593\(0 to 3);
              \$v6592\ := \$v6593\(4 to 35);
              case \$v6594\ is
              when "0001" =>
                \$15732\ := eclat_false;
              when "0000" =>
                \$15782_i\ := \$v6592\(0 to 31);
                \$15732\ := eclat_if(eclat_ge(\$15782_i\ & X"0000000" & X"0") & eclat_lt(\$15782_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v6591\ := \$15732\;
              if \$v6591\(0) = '1' then
                \$v6589\ := \$15724_len_aux3143361_arg\(0 to 35);
                \$v6590\ := \$v6589\(0 to 3);
                \$v6584\ := \$v6589\(4 to 35);
                case \$v6590\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$15772_forever3163360\;
                when "0000" =>
                  \$15780_i\ := \$v6584\(0 to 31);
                  \$v6588\ := \$$10696_ram_ptr_take\;
                  if \$v6588\(0) = '1' then
                    state_var7021 <= q_wait6587;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$15780_i\));
                    state_var7021 <= pause_getI6585;
                  end if;
                when others =>
                  
                end case;
              else
                \$15733\ := eclat_false;
                \$v6572\ := \$15733\;
                if \$v6572\(0) = '1' then
                  \$v6570\ := \$15724_len_aux3143361_arg\(0 to 35);
                  \$v6571\ := \$v6570\(0 to 3);
                  \$v6565\ := \$v6570\(4 to 35);
                  case \$v6571\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15746_forever3163359\;
                  when "0000" =>
                    \$15754_i\ := \$v6565\(0 to 31);
                    \$v6569\ := \$$10696_ram_ptr_take\;
                    if \$v6569\(0) = '1' then
                      state_var7021 <= q_wait6568;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15754_i\));
                      state_var7021 <= pause_getI6566;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15724_len_aux3143361_result\ := \$15724_len_aux3143361_arg\(36 to 67);
                  \$15622\ := \$15724_len_aux3143361_result\;
                  \$v6564\ := \$$10702_brk_ptr_take\;
                  if \$v6564\(0) = '1' then
                    state_var7021 <= q_wait6563;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6561;
                  end if;
                end if;
              end if;
            when \$15746_forever3163359\ =>
              state_var7021 <= \$15750_forever3163133\;
            when \$15750_forever3163133\ =>
              state_var7021 <= \$15750_forever3163133\;
            when \$15772_forever3163360\ =>
              state_var7021 <= \$15776_forever3163133\;
            when \$15776_forever3163133\ =>
              state_var7021 <= \$15776_forever3163133\;
            when \$15788_get_int268\ =>
              \$v6994\ := \$$10701_pos_ptr_take\;
              if \$v6994\(0) = '1' then
                state_var7021 <= q_wait6993;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6991;
              end if;
            when pause_getI3378 =>
              state_var7021 <= pause_getII3379;
            when pause_getI3397 =>
              state_var7021 <= pause_getII3398;
            when pause_getI3404 =>
              state_var7021 <= pause_getII3405;
            when pause_getI3418 =>
              state_var7021 <= pause_getII3419;
            when pause_getI3425 =>
              state_var7021 <= pause_getII3426;
            when pause_getI3433 =>
              state_var7021 <= pause_getII3434;
            when pause_getI3443 =>
              state_var7021 <= pause_getII3444;
            when pause_getI3450 =>
              state_var7021 <= pause_getII3451;
            when pause_getI3459 =>
              state_var7021 <= pause_getII3460;
            when pause_getI3471 =>
              state_var7021 <= pause_getII3472;
            when pause_getI3478 =>
              state_var7021 <= pause_getII3479;
            when pause_getI3487 =>
              state_var7021 <= pause_getII3488;
            when pause_getI3494 =>
              state_var7021 <= pause_getII3495;
            when pause_getI3505 =>
              state_var7021 <= pause_getII3506;
            when pause_getI3511 =>
              state_var7021 <= pause_getII3512;
            when pause_getI3519 =>
              state_var7021 <= pause_getII3520;
            when pause_getI3528 =>
              state_var7021 <= pause_getII3529;
            when pause_getI3536 =>
              state_var7021 <= pause_getII3537;
            when pause_getI3540 =>
              state_var7021 <= pause_getII3541;
            when pause_getI3548 =>
              state_var7021 <= pause_getII3549;
            when pause_getI3553 =>
              state_var7021 <= pause_getII3554;
            when pause_getI3557 =>
              state_var7021 <= pause_getII3558;
            when pause_getI3568 =>
              state_var7021 <= pause_getII3569;
            when pause_getI3572 =>
              state_var7021 <= pause_getII3573;
            when pause_getI3581 =>
              state_var7021 <= pause_getII3582;
            when pause_getI3587 =>
              state_var7021 <= pause_getII3588;
            when pause_getI3597 =>
              state_var7021 <= pause_getII3598;
            when pause_getI3605 =>
              state_var7021 <= pause_getII3606;
            when pause_getI3609 =>
              state_var7021 <= pause_getII3610;
            when pause_getI3617 =>
              state_var7021 <= pause_getII3618;
            when pause_getI3622 =>
              state_var7021 <= pause_getII3623;
            when pause_getI3626 =>
              state_var7021 <= pause_getII3627;
            when pause_getI3638 =>
              state_var7021 <= pause_getII3639;
            when pause_getI3644 =>
              state_var7021 <= pause_getII3645;
            when pause_getI3656 =>
              state_var7021 <= pause_getII3657;
            when pause_getI3668 =>
              state_var7021 <= pause_getII3669;
            when pause_getI3675 =>
              state_var7021 <= pause_getII3676;
            when pause_getI3684 =>
              state_var7021 <= pause_getII3685;
            when pause_getI3690 =>
              state_var7021 <= pause_getII3691;
            when pause_getI3695 =>
              state_var7021 <= pause_getII3696;
            when pause_getI3706 =>
              state_var7021 <= pause_getII3707;
            when pause_getI3712 =>
              state_var7021 <= pause_getII3713;
            when pause_getI3725 =>
              state_var7021 <= pause_getII3726;
            when pause_getI3733 =>
              state_var7021 <= pause_getII3734;
            when pause_getI3737 =>
              state_var7021 <= pause_getII3738;
            when pause_getI3741 =>
              state_var7021 <= pause_getII3742;
            when pause_getI3749 =>
              state_var7021 <= pause_getII3750;
            when pause_getI3754 =>
              state_var7021 <= pause_getII3755;
            when pause_getI3758 =>
              state_var7021 <= pause_getII3759;
            when pause_getI3762 =>
              state_var7021 <= pause_getII3763;
            when pause_getI3770 =>
              state_var7021 <= pause_getII3771;
            when pause_getI3778 =>
              state_var7021 <= pause_getII3779;
            when pause_getI3782 =>
              state_var7021 <= pause_getII3783;
            when pause_getI3790 =>
              state_var7021 <= pause_getII3791;
            when pause_getI3795 =>
              state_var7021 <= pause_getII3796;
            when pause_getI3799 =>
              state_var7021 <= pause_getII3800;
            when pause_getI3810 =>
              state_var7021 <= pause_getII3811;
            when pause_getI3814 =>
              state_var7021 <= pause_getII3815;
            when pause_getI3825 =>
              state_var7021 <= pause_getII3826;
            when pause_getI3829 =>
              state_var7021 <= pause_getII3830;
            when pause_getI3840 =>
              state_var7021 <= pause_getII3841;
            when pause_getI3844 =>
              state_var7021 <= pause_getII3845;
            when pause_getI3853 =>
              state_var7021 <= pause_getII3854;
            when pause_getI3861 =>
              state_var7021 <= pause_getII3862;
            when pause_getI3865 =>
              state_var7021 <= pause_getII3866;
            when pause_getI3869 =>
              state_var7021 <= pause_getII3870;
            when pause_getI3877 =>
              state_var7021 <= pause_getII3878;
            when pause_getI3882 =>
              state_var7021 <= pause_getII3883;
            when pause_getI3886 =>
              state_var7021 <= pause_getII3887;
            when pause_getI3897 =>
              state_var7021 <= pause_getII3898;
            when pause_getI3901 =>
              state_var7021 <= pause_getII3902;
            when pause_getI3912 =>
              state_var7021 <= pause_getII3913;
            when pause_getI3916 =>
              state_var7021 <= pause_getII3917;
            when pause_getI3925 =>
              state_var7021 <= pause_getII3926;
            when pause_getI3933 =>
              state_var7021 <= pause_getII3934;
            when pause_getI3937 =>
              state_var7021 <= pause_getII3938;
            when pause_getI3941 =>
              state_var7021 <= pause_getII3942;
            when pause_getI3949 =>
              state_var7021 <= pause_getII3950;
            when pause_getI3954 =>
              state_var7021 <= pause_getII3955;
            when pause_getI3958 =>
              state_var7021 <= pause_getII3959;
            when pause_getI3969 =>
              state_var7021 <= pause_getII3970;
            when pause_getI3973 =>
              state_var7021 <= pause_getII3974;
            when pause_getI3984 =>
              state_var7021 <= pause_getII3985;
            when pause_getI3988 =>
              state_var7021 <= pause_getII3989;
            when pause_getI3997 =>
              state_var7021 <= pause_getII3998;
            when pause_getI4005 =>
              state_var7021 <= pause_getII4006;
            when pause_getI4009 =>
              state_var7021 <= pause_getII4010;
            when pause_getI4013 =>
              state_var7021 <= pause_getII4014;
            when pause_getI4021 =>
              state_var7021 <= pause_getII4022;
            when pause_getI4026 =>
              state_var7021 <= pause_getII4027;
            when pause_getI4030 =>
              state_var7021 <= pause_getII4031;
            when pause_getI4034 =>
              state_var7021 <= pause_getII4035;
            when pause_getI4043 =>
              state_var7021 <= pause_getII4044;
            when pause_getI4051 =>
              state_var7021 <= pause_getII4052;
            when pause_getI4055 =>
              state_var7021 <= pause_getII4056;
            when pause_getI4063 =>
              state_var7021 <= pause_getII4064;
            when pause_getI4068 =>
              state_var7021 <= pause_getII4069;
            when pause_getI4072 =>
              state_var7021 <= pause_getII4073;
            when pause_getI4076 =>
              state_var7021 <= pause_getII4077;
            when pause_getI4081 =>
              state_var7021 <= pause_getII4082;
            when pause_getI4094 =>
              state_var7021 <= pause_getII4095;
            when pause_getI4098 =>
              state_var7021 <= pause_getII4099;
            when pause_getI4109 =>
              state_var7021 <= pause_getII4110;
            when pause_getI4117 =>
              state_var7021 <= pause_getII4118;
            when pause_getI4121 =>
              state_var7021 <= pause_getII4122;
            when pause_getI4125 =>
              state_var7021 <= pause_getII4126;
            when pause_getI4133 =>
              state_var7021 <= pause_getII4134;
            when pause_getI4138 =>
              state_var7021 <= pause_getII4139;
            when pause_getI4142 =>
              state_var7021 <= pause_getII4143;
            when pause_getI4156 =>
              state_var7021 <= pause_getII4157;
            when pause_getI4160 =>
              state_var7021 <= pause_getII4161;
            when pause_getI4169 =>
              state_var7021 <= pause_getII4170;
            when pause_getI4177 =>
              state_var7021 <= pause_getII4178;
            when pause_getI4181 =>
              state_var7021 <= pause_getII4182;
            when pause_getI4185 =>
              state_var7021 <= pause_getII4186;
            when pause_getI4193 =>
              state_var7021 <= pause_getII4194;
            when pause_getI4198 =>
              state_var7021 <= pause_getII4199;
            when pause_getI4202 =>
              state_var7021 <= pause_getII4203;
            when pause_getI4207 =>
              state_var7021 <= pause_getII4208;
            when pause_getI4220 =>
              state_var7021 <= pause_getII4221;
            when pause_getI4224 =>
              state_var7021 <= pause_getII4225;
            when pause_getI4233 =>
              state_var7021 <= pause_getII4234;
            when pause_getI4241 =>
              state_var7021 <= pause_getII4242;
            when pause_getI4245 =>
              state_var7021 <= pause_getII4246;
            when pause_getI4249 =>
              state_var7021 <= pause_getII4250;
            when pause_getI4257 =>
              state_var7021 <= pause_getII4258;
            when pause_getI4262 =>
              state_var7021 <= pause_getII4263;
            when pause_getI4266 =>
              state_var7021 <= pause_getII4267;
            when pause_getI4271 =>
              state_var7021 <= pause_getII4272;
            when pause_getI4284 =>
              state_var7021 <= pause_getII4285;
            when pause_getI4288 =>
              state_var7021 <= pause_getII4289;
            when pause_getI4297 =>
              state_var7021 <= pause_getII4298;
            when pause_getI4305 =>
              state_var7021 <= pause_getII4306;
            when pause_getI4309 =>
              state_var7021 <= pause_getII4310;
            when pause_getI4313 =>
              state_var7021 <= pause_getII4314;
            when pause_getI4321 =>
              state_var7021 <= pause_getII4322;
            when pause_getI4326 =>
              state_var7021 <= pause_getII4327;
            when pause_getI4330 =>
              state_var7021 <= pause_getII4331;
            when pause_getI4335 =>
              state_var7021 <= pause_getII4336;
            when pause_getI4348 =>
              state_var7021 <= pause_getII4349;
            when pause_getI4352 =>
              state_var7021 <= pause_getII4353;
            when pause_getI4361 =>
              state_var7021 <= pause_getII4362;
            when pause_getI4369 =>
              state_var7021 <= pause_getII4370;
            when pause_getI4373 =>
              state_var7021 <= pause_getII4374;
            when pause_getI4377 =>
              state_var7021 <= pause_getII4378;
            when pause_getI4385 =>
              state_var7021 <= pause_getII4386;
            when pause_getI4390 =>
              state_var7021 <= pause_getII4391;
            when pause_getI4394 =>
              state_var7021 <= pause_getII4395;
            when pause_getI4404 =>
              state_var7021 <= pause_getII4405;
            when pause_getI4411 =>
              state_var7021 <= pause_getII4412;
            when pause_getI4426 =>
              state_var7021 <= pause_getII4427;
            when pause_getI4430 =>
              state_var7021 <= pause_getII4431;
            when pause_getI4441 =>
              state_var7021 <= pause_getII4442;
            when pause_getI4445 =>
              state_var7021 <= pause_getII4446;
            when pause_getI4454 =>
              state_var7021 <= pause_getII4455;
            when pause_getI4462 =>
              state_var7021 <= pause_getII4463;
            when pause_getI4466 =>
              state_var7021 <= pause_getII4467;
            when pause_getI4470 =>
              state_var7021 <= pause_getII4471;
            when pause_getI4478 =>
              state_var7021 <= pause_getII4479;
            when pause_getI4483 =>
              state_var7021 <= pause_getII4484;
            when pause_getI4487 =>
              state_var7021 <= pause_getII4488;
            when pause_getI4497 =>
              state_var7021 <= pause_getII4498;
            when pause_getI4504 =>
              state_var7021 <= pause_getII4505;
            when pause_getI4519 =>
              state_var7021 <= pause_getII4520;
            when pause_getI4523 =>
              state_var7021 <= pause_getII4524;
            when pause_getI4534 =>
              state_var7021 <= pause_getII4535;
            when pause_getI4538 =>
              state_var7021 <= pause_getII4539;
            when pause_getI4547 =>
              state_var7021 <= pause_getII4548;
            when pause_getI4555 =>
              state_var7021 <= pause_getII4556;
            when pause_getI4559 =>
              state_var7021 <= pause_getII4560;
            when pause_getI4563 =>
              state_var7021 <= pause_getII4564;
            when pause_getI4571 =>
              state_var7021 <= pause_getII4572;
            when pause_getI4576 =>
              state_var7021 <= pause_getII4577;
            when pause_getI4580 =>
              state_var7021 <= pause_getII4581;
            when pause_getI4590 =>
              state_var7021 <= pause_getII4591;
            when pause_getI4597 =>
              state_var7021 <= pause_getII4598;
            when pause_getI4612 =>
              state_var7021 <= pause_getII4613;
            when pause_getI4616 =>
              state_var7021 <= pause_getII4617;
            when pause_getI4627 =>
              state_var7021 <= pause_getII4628;
            when pause_getI4631 =>
              state_var7021 <= pause_getII4632;
            when pause_getI4642 =>
              state_var7021 <= pause_getII4643;
            when pause_getI4650 =>
              state_var7021 <= pause_getII4651;
            when pause_getI4654 =>
              state_var7021 <= pause_getII4655;
            when pause_getI4658 =>
              state_var7021 <= pause_getII4659;
            when pause_getI4666 =>
              state_var7021 <= pause_getII4667;
            when pause_getI4671 =>
              state_var7021 <= pause_getII4672;
            when pause_getI4675 =>
              state_var7021 <= pause_getII4676;
            when pause_getI4714 =>
              state_var7021 <= pause_getII4715;
            when pause_getI4721 =>
              state_var7021 <= pause_getII4722;
            when pause_getI4738 =>
              state_var7021 <= pause_getII4739;
            when pause_getI4742 =>
              state_var7021 <= pause_getII4743;
            when pause_getI4753 =>
              state_var7021 <= pause_getII4754;
            when pause_getI4757 =>
              state_var7021 <= pause_getII4758;
            when pause_getI4766 =>
              state_var7021 <= pause_getII4767;
            when pause_getI4774 =>
              state_var7021 <= pause_getII4775;
            when pause_getI4778 =>
              state_var7021 <= pause_getII4779;
            when pause_getI4782 =>
              state_var7021 <= pause_getII4783;
            when pause_getI4790 =>
              state_var7021 <= pause_getII4791;
            when pause_getI4795 =>
              state_var7021 <= pause_getII4796;
            when pause_getI4799 =>
              state_var7021 <= pause_getII4800;
            when pause_getI4818 =>
              state_var7021 <= pause_getII4819;
            when pause_getI4822 =>
              state_var7021 <= pause_getII4823;
            when pause_getI4833 =>
              state_var7021 <= pause_getII4834;
            when pause_getI4837 =>
              state_var7021 <= pause_getII4838;
            when pause_getI4846 =>
              state_var7021 <= pause_getII4847;
            when pause_getI4854 =>
              state_var7021 <= pause_getII4855;
            when pause_getI4858 =>
              state_var7021 <= pause_getII4859;
            when pause_getI4862 =>
              state_var7021 <= pause_getII4863;
            when pause_getI4870 =>
              state_var7021 <= pause_getII4871;
            when pause_getI4875 =>
              state_var7021 <= pause_getII4876;
            when pause_getI4879 =>
              state_var7021 <= pause_getII4880;
            when pause_getI4897 =>
              state_var7021 <= pause_getII4898;
            when pause_getI4901 =>
              state_var7021 <= pause_getII4902;
            when pause_getI4912 =>
              state_var7021 <= pause_getII4913;
            when pause_getI4916 =>
              state_var7021 <= pause_getII4917;
            when pause_getI4925 =>
              state_var7021 <= pause_getII4926;
            when pause_getI4933 =>
              state_var7021 <= pause_getII4934;
            when pause_getI4937 =>
              state_var7021 <= pause_getII4938;
            when pause_getI4941 =>
              state_var7021 <= pause_getII4942;
            when pause_getI4949 =>
              state_var7021 <= pause_getII4950;
            when pause_getI4954 =>
              state_var7021 <= pause_getII4955;
            when pause_getI4958 =>
              state_var7021 <= pause_getII4959;
            when pause_getI4976 =>
              state_var7021 <= pause_getII4977;
            when pause_getI4980 =>
              state_var7021 <= pause_getII4981;
            when pause_getI4991 =>
              state_var7021 <= pause_getII4992;
            when pause_getI4995 =>
              state_var7021 <= pause_getII4996;
            when pause_getI5004 =>
              state_var7021 <= pause_getII5005;
            when pause_getI5012 =>
              state_var7021 <= pause_getII5013;
            when pause_getI5016 =>
              state_var7021 <= pause_getII5017;
            when pause_getI5020 =>
              state_var7021 <= pause_getII5021;
            when pause_getI5028 =>
              state_var7021 <= pause_getII5029;
            when pause_getI5033 =>
              state_var7021 <= pause_getII5034;
            when pause_getI5037 =>
              state_var7021 <= pause_getII5038;
            when pause_getI5055 =>
              state_var7021 <= pause_getII5056;
            when pause_getI5059 =>
              state_var7021 <= pause_getII5060;
            when pause_getI5070 =>
              state_var7021 <= pause_getII5071;
            when pause_getI5074 =>
              state_var7021 <= pause_getII5075;
            when pause_getI5083 =>
              state_var7021 <= pause_getII5084;
            when pause_getI5091 =>
              state_var7021 <= pause_getII5092;
            when pause_getI5095 =>
              state_var7021 <= pause_getII5096;
            when pause_getI5099 =>
              state_var7021 <= pause_getII5100;
            when pause_getI5107 =>
              state_var7021 <= pause_getII5108;
            when pause_getI5112 =>
              state_var7021 <= pause_getII5113;
            when pause_getI5116 =>
              state_var7021 <= pause_getII5117;
            when pause_getI5134 =>
              state_var7021 <= pause_getII5135;
            when pause_getI5138 =>
              state_var7021 <= pause_getII5139;
            when pause_getI5149 =>
              state_var7021 <= pause_getII5150;
            when pause_getI5153 =>
              state_var7021 <= pause_getII5154;
            when pause_getI5162 =>
              state_var7021 <= pause_getII5163;
            when pause_getI5170 =>
              state_var7021 <= pause_getII5171;
            when pause_getI5174 =>
              state_var7021 <= pause_getII5175;
            when pause_getI5178 =>
              state_var7021 <= pause_getII5179;
            when pause_getI5186 =>
              state_var7021 <= pause_getII5187;
            when pause_getI5191 =>
              state_var7021 <= pause_getII5192;
            when pause_getI5195 =>
              state_var7021 <= pause_getII5196;
            when pause_getI5204 =>
              state_var7021 <= pause_getII5205;
            when pause_getI5212 =>
              state_var7021 <= pause_getII5213;
            when pause_getI5216 =>
              state_var7021 <= pause_getII5217;
            when pause_getI5220 =>
              state_var7021 <= pause_getII5221;
            when pause_getI5228 =>
              state_var7021 <= pause_getII5229;
            when pause_getI5233 =>
              state_var7021 <= pause_getII5234;
            when pause_getI5237 =>
              state_var7021 <= pause_getII5238;
            when pause_getI5251 =>
              state_var7021 <= pause_getII5252;
            when pause_getI5255 =>
              state_var7021 <= pause_getII5256;
            when pause_getI5263 =>
              state_var7021 <= pause_getII5264;
            when pause_getI5271 =>
              state_var7021 <= pause_getII5272;
            when pause_getI5278 =>
              state_var7021 <= pause_getII5279;
            when pause_getI5285 =>
              state_var7021 <= pause_getII5286;
            when pause_getI5290 =>
              state_var7021 <= pause_getII5291;
            when pause_getI5299 =>
              state_var7021 <= pause_getII5300;
            when pause_getI5305 =>
              state_var7021 <= pause_getII5306;
            when pause_getI5310 =>
              state_var7021 <= pause_getII5311;
            when pause_getI5314 =>
              state_var7021 <= pause_getII5315;
            when pause_getI5326 =>
              state_var7021 <= pause_getII5327;
            when pause_getI5332 =>
              state_var7021 <= pause_getII5333;
            when pause_getI5343 =>
              state_var7021 <= pause_getII5344;
            when pause_getI5350 =>
              state_var7021 <= pause_getII5351;
            when pause_getI5359 =>
              state_var7021 <= pause_getII5360;
            when pause_getI5366 =>
              state_var7021 <= pause_getII5367;
            when pause_getI5376 =>
              state_var7021 <= pause_getII5377;
            when pause_getI5383 =>
              state_var7021 <= pause_getII5384;
            when pause_getI5400 =>
              state_var7021 <= pause_getII5401;
            when pause_getI5404 =>
              state_var7021 <= pause_getII5405;
            when pause_getI5416 =>
              state_var7021 <= pause_getII5417;
            when pause_getI5422 =>
              state_var7021 <= pause_getII5423;
            when pause_getI5431 =>
              state_var7021 <= pause_getII5432;
            when pause_getI5439 =>
              state_var7021 <= pause_getII5440;
            when pause_getI5443 =>
              state_var7021 <= pause_getII5444;
            when pause_getI5447 =>
              state_var7021 <= pause_getII5448;
            when pause_getI5455 =>
              state_var7021 <= pause_getII5456;
            when pause_getI5460 =>
              state_var7021 <= pause_getII5461;
            when pause_getI5464 =>
              state_var7021 <= pause_getII5465;
            when pause_getI5470 =>
              state_var7021 <= pause_getII5471;
            when pause_getI5477 =>
              state_var7021 <= pause_getII5478;
            when pause_getI5484 =>
              state_var7021 <= pause_getII5485;
            when pause_getI5489 =>
              state_var7021 <= pause_getII5490;
            when pause_getI5505 =>
              state_var7021 <= pause_getII5506;
            when pause_getI5511 =>
              state_var7021 <= pause_getII5512;
            when pause_getI5520 =>
              state_var7021 <= pause_getII5521;
            when pause_getI5528 =>
              state_var7021 <= pause_getII5529;
            when pause_getI5532 =>
              state_var7021 <= pause_getII5533;
            when pause_getI5536 =>
              state_var7021 <= pause_getII5537;
            when pause_getI5544 =>
              state_var7021 <= pause_getII5545;
            when pause_getI5549 =>
              state_var7021 <= pause_getII5550;
            when pause_getI5553 =>
              state_var7021 <= pause_getII5554;
            when pause_getI5565 =>
              state_var7021 <= pause_getII5566;
            when pause_getI5571 =>
              state_var7021 <= pause_getII5572;
            when pause_getI5601 =>
              state_var7021 <= pause_getII5602;
            when pause_getI5605 =>
              state_var7021 <= pause_getII5606;
            when pause_getI5613 =>
              state_var7021 <= pause_getII5614;
            when pause_getI5619 =>
              state_var7021 <= pause_getII5620;
            when pause_getI5640 =>
              state_var7021 <= pause_getII5641;
            when pause_getI5644 =>
              state_var7021 <= pause_getII5645;
            when pause_getI5652 =>
              state_var7021 <= pause_getII5653;
            when pause_getI5657 =>
              state_var7021 <= pause_getII5658;
            when pause_getI5661 =>
              state_var7021 <= pause_getII5662;
            when pause_getI5665 =>
              state_var7021 <= pause_getII5666;
            when pause_getI5669 =>
              state_var7021 <= pause_getII5670;
            when pause_getI5677 =>
              state_var7021 <= pause_getII5678;
            when pause_getI5682 =>
              state_var7021 <= pause_getII5683;
            when pause_getI5686 =>
              state_var7021 <= pause_getII5687;
            when pause_getI5698 =>
              state_var7021 <= pause_getII5699;
            when pause_getI5704 =>
              state_var7021 <= pause_getII5705;
            when pause_getI5715 =>
              state_var7021 <= pause_getII5716;
            when pause_getI5722 =>
              state_var7021 <= pause_getII5723;
            when pause_getI5731 =>
              state_var7021 <= pause_getII5732;
            when pause_getI5737 =>
              state_var7021 <= pause_getII5738;
            when pause_getI5749 =>
              state_var7021 <= pause_getII5750;
            when pause_getI5755 =>
              state_var7021 <= pause_getII5756;
            when pause_getI5766 =>
              state_var7021 <= pause_getII5767;
            when pause_getI5773 =>
              state_var7021 <= pause_getII5774;
            when pause_getI5782 =>
              state_var7021 <= pause_getII5783;
            when pause_getI5788 =>
              state_var7021 <= pause_getII5789;
            when pause_getI5800 =>
              state_var7021 <= pause_getII5801;
            when pause_getI5806 =>
              state_var7021 <= pause_getII5807;
            when pause_getI5817 =>
              state_var7021 <= pause_getII5818;
            when pause_getI5824 =>
              state_var7021 <= pause_getII5825;
            when pause_getI5833 =>
              state_var7021 <= pause_getII5834;
            when pause_getI5839 =>
              state_var7021 <= pause_getII5840;
            when pause_getI5851 =>
              state_var7021 <= pause_getII5852;
            when pause_getI5857 =>
              state_var7021 <= pause_getII5858;
            when pause_getI5867 =>
              state_var7021 <= pause_getII5868;
            when pause_getI5874 =>
              state_var7021 <= pause_getII5875;
            when pause_getI5883 =>
              state_var7021 <= pause_getII5884;
            when pause_getI5889 =>
              state_var7021 <= pause_getII5890;
            when pause_getI5893 =>
              state_var7021 <= pause_getII5894;
            when pause_getI5903 =>
              state_var7021 <= pause_getII5904;
            when pause_getI5911 =>
              state_var7021 <= pause_getII5912;
            when pause_getI5915 =>
              state_var7021 <= pause_getII5916;
            when pause_getI5923 =>
              state_var7021 <= pause_getII5924;
            when pause_getI5928 =>
              state_var7021 <= pause_getII5929;
            when pause_getI5932 =>
              state_var7021 <= pause_getII5933;
            when pause_getI5936 =>
              state_var7021 <= pause_getII5937;
            when pause_getI5948 =>
              state_var7021 <= pause_getII5949;
            when pause_getI5955 =>
              state_var7021 <= pause_getII5956;
            when pause_getI5961 =>
              state_var7021 <= pause_getII5962;
            when pause_getI5971 =>
              state_var7021 <= pause_getII5972;
            when pause_getI5978 =>
              state_var7021 <= pause_getII5979;
            when pause_getI5986 =>
              state_var7021 <= pause_getII5987;
            when pause_getI5995 =>
              state_var7021 <= pause_getII5996;
            when pause_getI6003 =>
              state_var7021 <= pause_getII6004;
            when pause_getI6007 =>
              state_var7021 <= pause_getII6008;
            when pause_getI6015 =>
              state_var7021 <= pause_getII6016;
            when pause_getI6020 =>
              state_var7021 <= pause_getII6021;
            when pause_getI6024 =>
              state_var7021 <= pause_getII6025;
            when pause_getI6029 =>
              state_var7021 <= pause_getII6030;
            when pause_getI6035 =>
              state_var7021 <= pause_getII6036;
            when pause_getI6046 =>
              state_var7021 <= pause_getII6047;
            when pause_getI6050 =>
              state_var7021 <= pause_getII6051;
            when pause_getI6060 =>
              state_var7021 <= pause_getII6061;
            when pause_getI6067 =>
              state_var7021 <= pause_getII6068;
            when pause_getI6075 =>
              state_var7021 <= pause_getII6076;
            when pause_getI6084 =>
              state_var7021 <= pause_getII6085;
            when pause_getI6092 =>
              state_var7021 <= pause_getII6093;
            when pause_getI6096 =>
              state_var7021 <= pause_getII6097;
            when pause_getI6104 =>
              state_var7021 <= pause_getII6105;
            when pause_getI6109 =>
              state_var7021 <= pause_getII6110;
            when pause_getI6113 =>
              state_var7021 <= pause_getII6114;
            when pause_getI6118 =>
              state_var7021 <= pause_getII6119;
            when pause_getI6124 =>
              state_var7021 <= pause_getII6125;
            when pause_getI6132 =>
              state_var7021 <= pause_getII6133;
            when pause_getI6136 =>
              state_var7021 <= pause_getII6137;
            when pause_getI6146 =>
              state_var7021 <= pause_getII6147;
            when pause_getI6154 =>
              state_var7021 <= pause_getII6155;
            when pause_getI6158 =>
              state_var7021 <= pause_getII6159;
            when pause_getI6166 =>
              state_var7021 <= pause_getII6167;
            when pause_getI6171 =>
              state_var7021 <= pause_getII6172;
            when pause_getI6175 =>
              state_var7021 <= pause_getII6176;
            when pause_getI6179 =>
              state_var7021 <= pause_getII6180;
            when pause_getI6188 =>
              state_var7021 <= pause_getII6189;
            when pause_getI6196 =>
              state_var7021 <= pause_getII6197;
            when pause_getI6200 =>
              state_var7021 <= pause_getII6201;
            when pause_getI6208 =>
              state_var7021 <= pause_getII6209;
            when pause_getI6213 =>
              state_var7021 <= pause_getII6214;
            when pause_getI6217 =>
              state_var7021 <= pause_getII6218;
            when pause_getI6228 =>
              state_var7021 <= pause_getII6229;
            when pause_getI6232 =>
              state_var7021 <= pause_getII6233;
            when pause_getI6242 =>
              state_var7021 <= pause_getII6243;
            when pause_getI6249 =>
              state_var7021 <= pause_getII6250;
            when pause_getI6257 =>
              state_var7021 <= pause_getII6258;
            when pause_getI6266 =>
              state_var7021 <= pause_getII6267;
            when pause_getI6274 =>
              state_var7021 <= pause_getII6275;
            when pause_getI6278 =>
              state_var7021 <= pause_getII6279;
            when pause_getI6286 =>
              state_var7021 <= pause_getII6287;
            when pause_getI6291 =>
              state_var7021 <= pause_getII6292;
            when pause_getI6295 =>
              state_var7021 <= pause_getII6296;
            when pause_getI6300 =>
              state_var7021 <= pause_getII6301;
            when pause_getI6306 =>
              state_var7021 <= pause_getII6307;
            when pause_getI6312 =>
              state_var7021 <= pause_getII6313;
            when pause_getI6319 =>
              state_var7021 <= pause_getII6320;
            when pause_getI6326 =>
              state_var7021 <= pause_getII6327;
            when pause_getI6337 =>
              state_var7021 <= pause_getII6338;
            when pause_getI6341 =>
              state_var7021 <= pause_getII6342;
            when pause_getI6346 =>
              state_var7021 <= pause_getII6347;
            when pause_getI6353 =>
              state_var7021 <= pause_getII6354;
            when pause_getI6360 =>
              state_var7021 <= pause_getII6361;
            when pause_getI6369 =>
              state_var7021 <= pause_getII6370;
            when pause_getI6373 =>
              state_var7021 <= pause_getII6374;
            when pause_getI6385 =>
              state_var7021 <= pause_getII6386;
            when pause_getI6393 =>
              state_var7021 <= pause_getII6394;
            when pause_getI6397 =>
              state_var7021 <= pause_getII6398;
            when pause_getI6401 =>
              state_var7021 <= pause_getII6402;
            when pause_getI6409 =>
              state_var7021 <= pause_getII6410;
            when pause_getI6414 =>
              state_var7021 <= pause_getII6415;
            when pause_getI6418 =>
              state_var7021 <= pause_getII6419;
            when pause_getI6429 =>
              state_var7021 <= pause_getII6430;
            when pause_getI6433 =>
              state_var7021 <= pause_getII6434;
            when pause_getI6437 =>
              state_var7021 <= pause_getII6438;
            when pause_getI6446 =>
              state_var7021 <= pause_getII6447;
            when pause_getI6454 =>
              state_var7021 <= pause_getII6455;
            when pause_getI6458 =>
              state_var7021 <= pause_getII6459;
            when pause_getI6466 =>
              state_var7021 <= pause_getII6467;
            when pause_getI6471 =>
              state_var7021 <= pause_getII6472;
            when pause_getI6475 =>
              state_var7021 <= pause_getII6476;
            when pause_getI6479 =>
              state_var7021 <= pause_getII6480;
            when pause_getI6489 =>
              state_var7021 <= pause_getII6490;
            when pause_getI6497 =>
              state_var7021 <= pause_getII6498;
            when pause_getI6501 =>
              state_var7021 <= pause_getII6502;
            when pause_getI6509 =>
              state_var7021 <= pause_getII6510;
            when pause_getI6514 =>
              state_var7021 <= pause_getII6515;
            when pause_getI6518 =>
              state_var7021 <= pause_getII6519;
            when pause_getI6522 =>
              state_var7021 <= pause_getII6523;
            when pause_getI6532 =>
              state_var7021 <= pause_getII6533;
            when pause_getI6540 =>
              state_var7021 <= pause_getII6541;
            when pause_getI6544 =>
              state_var7021 <= pause_getII6545;
            when pause_getI6552 =>
              state_var7021 <= pause_getII6553;
            when pause_getI6557 =>
              state_var7021 <= pause_getII6558;
            when pause_getI6561 =>
              state_var7021 <= pause_getII6562;
            when pause_getI6566 =>
              state_var7021 <= pause_getII6567;
            when pause_getI6585 =>
              state_var7021 <= pause_getII6586;
            when pause_getI6596 =>
              state_var7021 <= pause_getII6597;
            when pause_getI6601 =>
              state_var7021 <= pause_getII6602;
            when pause_getI6610 =>
              state_var7021 <= pause_getII6611;
            when pause_getI6618 =>
              state_var7021 <= pause_getII6619;
            when pause_getI6622 =>
              state_var7021 <= pause_getII6623;
            when pause_getI6630 =>
              state_var7021 <= pause_getII6631;
            when pause_getI6635 =>
              state_var7021 <= pause_getII6636;
            when pause_getI6639 =>
              state_var7021 <= pause_getII6640;
            when pause_getI6643 =>
              state_var7021 <= pause_getII6644;
            when pause_getI6653 =>
              state_var7021 <= pause_getII6654;
            when pause_getI6661 =>
              state_var7021 <= pause_getII6662;
            when pause_getI6665 =>
              state_var7021 <= pause_getII6666;
            when pause_getI6673 =>
              state_var7021 <= pause_getII6674;
            when pause_getI6678 =>
              state_var7021 <= pause_getII6679;
            when pause_getI6682 =>
              state_var7021 <= pause_getII6683;
            when pause_getI6686 =>
              state_var7021 <= pause_getII6687;
            when pause_getI6695 =>
              state_var7021 <= pause_getII6696;
            when pause_getI6703 =>
              state_var7021 <= pause_getII6704;
            when pause_getI6707 =>
              state_var7021 <= pause_getII6708;
            when pause_getI6715 =>
              state_var7021 <= pause_getII6716;
            when pause_getI6720 =>
              state_var7021 <= pause_getII6721;
            when pause_getI6724 =>
              state_var7021 <= pause_getII6725;
            when pause_getI6729 =>
              state_var7021 <= pause_getII6730;
            when pause_getI6748 =>
              state_var7021 <= pause_getII6749;
            when pause_getI6758 =>
              state_var7021 <= pause_getII6759;
            when pause_getI6762 =>
              state_var7021 <= pause_getII6763;
            when pause_getI6771 =>
              state_var7021 <= pause_getII6772;
            when pause_getI6779 =>
              state_var7021 <= pause_getII6780;
            when pause_getI6783 =>
              state_var7021 <= pause_getII6784;
            when pause_getI6791 =>
              state_var7021 <= pause_getII6792;
            when pause_getI6796 =>
              state_var7021 <= pause_getII6797;
            when pause_getI6800 =>
              state_var7021 <= pause_getII6801;
            when pause_getI6804 =>
              state_var7021 <= pause_getII6805;
            when pause_getI6814 =>
              state_var7021 <= pause_getII6815;
            when pause_getI6822 =>
              state_var7021 <= pause_getII6823;
            when pause_getI6826 =>
              state_var7021 <= pause_getII6827;
            when pause_getI6834 =>
              state_var7021 <= pause_getII6835;
            when pause_getI6839 =>
              state_var7021 <= pause_getII6840;
            when pause_getI6843 =>
              state_var7021 <= pause_getII6844;
            when pause_getI6847 =>
              state_var7021 <= pause_getII6848;
            when pause_getI6856 =>
              state_var7021 <= pause_getII6857;
            when pause_getI6864 =>
              state_var7021 <= pause_getII6865;
            when pause_getI6868 =>
              state_var7021 <= pause_getII6869;
            when pause_getI6876 =>
              state_var7021 <= pause_getII6877;
            when pause_getI6881 =>
              state_var7021 <= pause_getII6882;
            when pause_getI6885 =>
              state_var7021 <= pause_getII6886;
            when pause_getI6890 =>
              state_var7021 <= pause_getII6891;
            when pause_getI6909 =>
              state_var7021 <= pause_getII6910;
            when pause_getI6919 =>
              state_var7021 <= pause_getII6920;
            when pause_getI6923 =>
              state_var7021 <= pause_getII6924;
            when pause_getI6933 =>
              state_var7021 <= pause_getII6934;
            when pause_getI6941 =>
              state_var7021 <= pause_getII6942;
            when pause_getI6945 =>
              state_var7021 <= pause_getII6946;
            when pause_getI6953 =>
              state_var7021 <= pause_getII6954;
            when pause_getI6958 =>
              state_var7021 <= pause_getII6959;
            when pause_getI6962 =>
              state_var7021 <= pause_getII6963;
            when pause_getI6972 =>
              state_var7021 <= pause_getII6973;
            when pause_getI6976 =>
              state_var7021 <= pause_getII6977;
            when pause_getI6987 =>
              state_var7021 <= pause_getII6988;
            when pause_getI6991 =>
              state_var7021 <= pause_getII6992;
            when pause_getII3379 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10848\ := \$$10696_ram_value\;
              \$v3375\ := \$10848\(72 to 107);
              \$v3376\ := \$v3375\(0 to 3);
              \$v3374\ := \$v3375\(4 to 35);
              case \$v3376\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10859_forever3163136\;
              when "0000" =>
                \$10867_i\ := \$v3374\(0 to 31);
                \$10853\ := \$10867_i\;
                \$v3373\ := \$$10700_pc_ptr_take\;
                if \$v3373\(0) = '1' then
                  state_var7021 <= q_wait3372;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr_write\ <= 0;
                  \$$10700_pc_write_request\ <= '1';
                  \$$10700_pc_write\ <= \$10853\;
                  state_var7021 <= pause_setI3370;
                end if;
              when others =>
                
              end case;
            when pause_getII3398 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11100\ := \$$10696_ram_value\;
              \$v3395\ := \$$10696_ram_ptr_take\;
              if \$v3395\(0) = '1' then
                state_var7021 <= q_wait3394;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11098_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11099\(0 to 35) & \$11100\(36 to 71) & \$10814\(72 to 107);
                state_var7021 <= pause_setI3392;
              end if;
            when pause_getII3405 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11099\ := \$$10696_ram_value\;
              \$v3401\ := \$10828_c2_rib\;
              \$v3402\ := \$v3401\(0 to 3);
              \$v3396\ := \$v3401\(4 to 35);
              case \$v3402\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11113_forever3163151\;
              when "0000" =>
                \$11121_i\ := \$v3396\(0 to 31);
                \$v3400\ := \$$10696_ram_ptr_take\;
                if \$v3400\(0) = '1' then
                  state_var7021 <= q_wait3399;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11121_i\));
                  state_var7021 <= pause_getI3397;
                end if;
              when others =>
                
              end case;
            when pause_getII3419 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11149\ := \$$10696_ram_value\;
              \$v3416\ := \$$10696_ram_ptr_take\;
              if \$v3416\(0) = '1' then
                state_var7021 <= q_wait3415;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11147_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$11084\ & \$11148\(36 to 71) & \$11149\(72 to 107);
                state_var7021 <= pause_setI3413;
              end if;
            when pause_getII3426 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11148\ := \$$10696_ram_value\;
              \$v3422\ := \$10828_c2_rib\;
              \$v3423\ := \$v3422\(0 to 3);
              \$v3417\ := \$v3422\(4 to 35);
              case \$v3423\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11164_forever3163154\;
              when "0000" =>
                \$11172_i\ := \$v3417\(0 to 31);
                \$v3421\ := \$$10696_ram_ptr_take\;
                if \$v3421\(0) = '1' then
                  state_var7021 <= q_wait3420;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11172_i\));
                  state_var7021 <= pause_getI3418;
                end if;
              when others =>
                
              end case;
            when pause_getII3434 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11084\ := \$$10697_stack_value\;
              \$v3431\ := \$10828_c2_rib\;
              \$v3432\ := \$v3431\(0 to 3);
              \$v3412\ := \$v3431\(4 to 35);
              case \$v3432\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11139_forever3163153\;
              when "0000" =>
                \$11147_i\ := \$v3412\(0 to 31);
                \$v3429\ := \$10828_c2_rib\;
                \$v3430\ := \$v3429\(0 to 3);
                \$v3424\ := \$v3429\(4 to 35);
                case \$v3430\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$11177_forever3163155\;
                when "0000" =>
                  \$11185_i\ := \$v3424\(0 to 31);
                  \$v3428\ := \$$10696_ram_ptr_take\;
                  if \$v3428\(0) = '1' then
                    state_var7021 <= q_wait3427;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$11185_i\));
                    state_var7021 <= pause_getI3425;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII3444 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10915\ := \$$10696_ram_value\;
              \$v3441\ := \$$10696_ram_ptr_take\;
              if \$v3441\(0) = '1' then
                state_var7021 <= q_wait3440;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10913_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$10914\(0 to 35) & \$10915\(36 to 71) & \$10900\(72 to 107);
                state_var7021 <= pause_setI3438;
              end if;
            when pause_getII3451 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10914\ := \$$10696_ram_value\;
              \$v3447\ := \$10828_c2_rib\;
              \$v3448\ := \$v3447\(0 to 3);
              \$v3442\ := \$v3447\(4 to 35);
              case \$v3448\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10932_forever3163140\;
              when "0000" =>
                \$10940_i\ := \$v3442\(0 to 31);
                \$v3446\ := \$$10696_ram_ptr_take\;
                if \$v3446\(0) = '1' then
                  state_var7021 <= q_wait3445;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$10940_i\));
                  state_var7021 <= pause_getI3443;
                end if;
              when others =>
                
              end case;
            when pause_getII3460 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10900\ := \$$10696_ram_value\;
              \$v3456\ := \$10828_c2_rib\;
              \$v3457\ := \$v3456\(0 to 3);
              \$v3437\ := \$v3456\(4 to 35);
              case \$v3457\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field2_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10905_forever3163139\;
              when "0000" =>
                \$10913_i\ := \$v3437\(0 to 31);
                \$v3454\ := \$10828_c2_rib\;
                \$v3455\ := \$v3454\(0 to 3);
                \$v3449\ := \$v3454\(4 to 35);
                case \$v3455\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$10945_forever3163141\;
                when "0000" =>
                  \$10953_i\ := \$v3449\(0 to 31);
                  \$v3453\ := \$$10696_ram_ptr_take\;
                  if \$v3453\(0) = '1' then
                    state_var7021 <= q_wait3452;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$10953_i\));
                    state_var7021 <= pause_getI3450;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII3472 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10981\ := \$$10696_ram_value\;
              \$v3469\ := \$$10696_ram_ptr_take\;
              if \$v3469\(0) = '1' then
                state_var7021 <= q_wait3468;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10979_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$10898\(0 to 35) & \$10980\(36 to 71) & \$10981\(72 to 107);
                state_var7021 <= pause_setI3466;
              end if;
            when pause_getII3479 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10980\ := \$$10696_ram_value\;
              \$v3475\ := \$10828_c2_rib\;
              \$v3476\ := \$v3475\(0 to 3);
              \$v3470\ := \$v3475\(4 to 35);
              case \$v3476\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10998_forever3163144\;
              when "0000" =>
                \$11006_i\ := \$v3470\(0 to 31);
                \$v3474\ := \$$10696_ram_ptr_take\;
                if \$v3474\(0) = '1' then
                  state_var7021 <= q_wait3473;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11006_i\));
                  state_var7021 <= pause_getI3471;
                end if;
              when others =>
                
              end case;
            when pause_getII3488 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10898\ := \$$10696_ram_value\;
              \$v3484\ := \$10828_c2_rib\;
              \$v3485\ := \$v3484\(0 to 3);
              \$v3465\ := \$v3484\(4 to 35);
              case \$v3485\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10971_forever3163143\;
              when "0000" =>
                \$10979_i\ := \$v3465\(0 to 31);
                \$v3482\ := \$10828_c2_rib\;
                \$v3483\ := \$v3482\(0 to 3);
                \$v3477\ := \$v3482\(4 to 35);
                case \$v3483\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$11011_forever3163145\;
                when "0000" =>
                  \$11019_i\ := \$v3477\(0 to 31);
                  \$v3481\ := \$$10696_ram_ptr_take\;
                  if \$v3481\(0) = '1' then
                    state_var7021 <= q_wait3480;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$11019_i\));
                    state_var7021 <= pause_getI3478;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII3495 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11048\ := \$$10696_ram_value\;
              \$11036_loop3073149_arg\ := \$11048\(36 to 71) & eclat_unit;
              state_var7021 <= \$11036_loop3073149\;
            when pause_getII3506 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11042\ := \$$10696_ram_value\;
              \$v3502\ := \$11042\(72 to 107);
              \$v3503\ := \$v3502\(0 to 3);
              \$v3501\ := \$v3502\(4 to 35);
              case \$v3503\ is
              when "0001" =>
                \$11047\ := eclat_false;
              when "0000" =>
                \$11067_i\ := \$v3501\(0 to 31);
                \$11047\ := eclat_if(eclat_ge(\$11067_i\ & X"0000000" & X"0") & eclat_lt(\$11067_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3500\ := \$11047\;
              if \$v3500\(0) = '1' then
                \$11036_loop3073149_result\ := \$11036_loop3073149_arg\(0 to 35);
                \$10897_k\ := \$11036_loop3073149_result\;
                \$v3491\ := \$10897_k\;
                \$v3492\ := \$v3491\(0 to 3);
                \$v3486\ := \$v3491\(4 to 35);
                case \$v3492\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$11024_forever3163146\;
                when "0000" =>
                  \$11032_i\ := \$v3486\(0 to 31);
                  \$v3490\ := \$$10696_ram_ptr_take\;
                  if \$v3490\(0) = '1' then
                    state_var7021 <= q_wait3489;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$11032_i\));
                    state_var7021 <= pause_getI3487;
                  end if;
                when others =>
                  
                end case;
              else
                \$v3498\ := \$11036_loop3073149_arg\(0 to 35);
                \$v3499\ := \$v3498\(0 to 3);
                \$v3493\ := \$v3498\(4 to 35);
                case \$v3499\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$11057_forever3163147\;
                when "0000" =>
                  \$11065_i\ := \$v3493\(0 to 31);
                  \$v3497\ := \$$10696_ram_ptr_take\;
                  if \$v3497\(0) = '1' then
                    state_var7021 <= q_wait3496;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$11065_i\));
                    state_var7021 <= pause_getI3494;
                  end if;
                when others =>
                  
                end case;
              end if;
            when pause_getII3512 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$10896\ := \$$10697_stack_value\;
              \$11036_loop3073149_arg\ := "0000" & \$10896\ & eclat_unit;
              state_var7021 <= \$11036_loop3073149\;
            when pause_getII3520 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$11232\ := \$$10698_heap_value\;
              \$11223\ := "0000" & \$11232\;
              \$11196_loop2913158_arg\ := eclat_sub(\$11196_loop2913158_arg\(0 to 31) & X"0000000" & X"1") & \$11223\ & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var7021 <= \$11196_loop2913158\;
            when pause_getII3529 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$11230\ := \$$10698_heap_value\;
              \$v3527\ := \$$10696_ram_ptr_take\;
              if \$v3527\(0) = '1' then
                state_var7021 <= q_wait3526;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3523\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11230\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11219\ & \$11196_loop2913158_arg\(32 to 67) & "0001" & \$v3523\;
                state_var7021 <= pause_setI3524;
              end if;
            when pause_getII3537 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11228_i\ := \$$10702_brk_value\;
              \$v3535\ := \$$10698_heap_ptr_take\;
              if \$v3535\(0) = '1' then
                state_var7021 <= q_wait3534;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11228_i\;
                state_var7021 <= pause_setI3532;
              end if;
            when pause_getII3541 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11228_i\ := \$$10702_brk_value\;
              \$v3535\ := \$$10698_heap_ptr_take\;
              if \$v3535\(0) = '1' then
                state_var7021 <= q_wait3534;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11228_i\;
                state_var7021 <= pause_setI3532;
              end if;
            when pause_getII3549 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11236\ := \$$10702_brk_value\;
              \$v3547\ := \$$10702_brk_ptr_take\;
              if \$v3547\(0) = '1' then
                state_var7021 <= q_wait3546;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11236\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3544;
              end if;
            when pause_getII3554 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11222\ := \$$10695_limit_value\;
              \$v3552\ := eclat_eq(\$11221\ & eclat_sub(\$11222\ & X"0000000" & X"1"));
              if \$v3552\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11244_forever3163156\;
              else
                \$v3551\ := \$$10702_brk_ptr_take\;
                if \$v3551\(0) = '1' then
                  state_var7021 <= q_wait3550;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI3548;
                end if;
              end if;
            when pause_getII3558 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11221\ := \$$10702_brk_value\;
              \$v3556\ := \$$10695_limit_ptr_take\;
              if \$v3556\(0) = '1' then
                state_var7021 <= q_wait3555;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3553;
              end if;
            when pause_getII3569 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11214\ := \$$10696_ram_value\;
              \$v3566\ := \$11214\(36 to 71);
              \$v3567\ := \$v3566\(0 to 3);
              \$v3565\ := \$v3566\(4 to 35);
              case \$v3567\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11259_forever3163157\;
              when "0000" =>
                \$11267_i\ := \$v3565\(0 to 31);
                \$11218\ := \$11267_i\;
                \$v3564\ := \$$10697_stack_ptr_take\;
                if \$v3564\(0) = '1' then
                  state_var7021 <= q_wait3563;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11218\;
                  state_var7021 <= pause_setI3561;
                end if;
              when others =>
                
              end case;
            when pause_getII3573 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11213\ := \$$10697_stack_value\;
              \$v3571\ := \$$10696_ram_ptr_take\;
              if \$v3571\(0) = '1' then
                state_var7021 <= q_wait3570;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11213\));
                state_var7021 <= pause_getI3568;
              end if;
            when pause_getII3582 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10833\ := \$$10696_ram_value\;
              \$v3578\ := \$10833\(0 to 35);
              \$v3579\ := \$v3578\(0 to 3);
              \$v3577\ := \$v3578\(4 to 35);
              case \$v3579\ is
              when "0000" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't inf_of_Int"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11272_forever3163159\;
              when "0001" =>
                \$11280_i\ := \$v3577\(0 to 31);
                \$10838_nargs\ := \$11280_i\;
                \$11196_loop2913158_arg\ := \$10838_nargs\ & \$10828_c2_rib\ & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
                state_var7021 <= \$11196_loop2913158\;
              when others =>
                
              end case;
            when pause_getII3588 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$11298\ := \$$10698_heap_value\;
              \$10828_c2_rib\ := "0000" & \$11298\;
              \$v3585\ := \$10819\(0 to 35);
              \$v3586\ := \$v3585\(0 to 3);
              \$v3580\ := \$v3585\(4 to 35);
              case \$v3586\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11285_forever3163160\;
              when "0000" =>
                \$11293_i\ := \$v3580\(0 to 31);
                \$v3584\ := \$$10696_ram_ptr_take\;
                if \$v3584\(0) = '1' then
                  state_var7021 <= q_wait3583;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11293_i\));
                  state_var7021 <= pause_getI3581;
                end if;
              when others =>
                
              end case;
            when pause_getII3598 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$11296\ := \$$10698_heap_value\;
              \$v3596\ := \$$10696_ram_ptr_take\;
              if \$v3596\(0) = '1' then
                state_var7021 <= q_wait3595;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3591\ := X"0000000" & X"0";
                \$v3592\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11296\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v3591\ & \$10818_proc\ & "0001" & \$v3592\;
                state_var7021 <= pause_setI3593;
              end if;
            when pause_getII3606 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11294_i\ := \$$10702_brk_value\;
              \$v3604\ := \$$10698_heap_ptr_take\;
              if \$v3604\(0) = '1' then
                state_var7021 <= q_wait3603;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11294_i\;
                state_var7021 <= pause_setI3601;
              end if;
            when pause_getII3610 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11294_i\ := \$$10702_brk_value\;
              \$v3604\ := \$$10698_heap_ptr_take\;
              if \$v3604\(0) = '1' then
                state_var7021 <= q_wait3603;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11294_i\;
                state_var7021 <= pause_setI3601;
              end if;
            when pause_getII3618 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11303\ := \$$10702_brk_value\;
              \$v3616\ := \$$10702_brk_ptr_take\;
              if \$v3616\(0) = '1' then
                state_var7021 <= q_wait3615;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11303\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3613;
              end if;
            when pause_getII3623 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$10827\ := \$$10695_limit_value\;
              \$v3621\ := eclat_eq(\$10826\ & eclat_sub(\$10827\ & X"0000000" & X"1"));
              if \$v3621\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11311_forever3163161\;
              else
                \$v3620\ := \$$10702_brk_ptr_take\;
                if \$v3620\(0) = '1' then
                  state_var7021 <= q_wait3619;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI3617;
                end if;
              end if;
            when pause_getII3627 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10826\ := \$$10702_brk_value\;
              \$v3625\ := \$$10695_limit_ptr_take\;
              if \$v3625\(0) = '1' then
                state_var7021 <= q_wait3624;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3622;
              end if;
            when pause_getII3639 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11486\ := \$$10696_ram_value\;
              \$v3635\ := \$11486\(72 to 107);
              \$v3636\ := \$v3635\(0 to 3);
              \$v3634\ := \$v3635\(4 to 35);
              case \$v3636\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11496_forever3163171\;
              when "0000" =>
                \$11504_i\ := \$v3634\(0 to 31);
                \$11491\ := \$11504_i\;
                \$v3633\ := \$$10700_pc_ptr_take\;
                if \$v3633\(0) = '1' then
                  state_var7021 <= q_wait3632;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr_write\ <= 0;
                  \$$10700_pc_write_request\ <= '1';
                  \$$10700_pc_write\ <= \$11491\;
                  state_var7021 <= pause_setI3630;
                end if;
              when others =>
                
              end case;
            when pause_getII3645 =>
              \$$10700_pc_ptr_take\(0) := '0';
              \$11485\ := \$$10700_pc_value\;
              \$v3642\ := "0000" & \$11485\;
              \$v3643\ := \$v3642\(0 to 3);
              \$v3637\ := \$v3642\(4 to 35);
              case \$v3643\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11510_forever3163172\;
              when "0000" =>
                \$11518_i\ := \$v3637\(0 to 31);
                \$v3641\ := \$$10696_ram_ptr_take\;
                if \$v3641\(0) = '1' then
                  state_var7021 <= q_wait3640;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11518_i\));
                  state_var7021 <= pause_getI3638;
                end if;
              when others =>
                
              end case;
            when pause_getII3657 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11333\ := \$$10696_ram_value\;
              \$v3653\ := \$11333\(72 to 107);
              \$v3654\ := \$v3653\(0 to 3);
              \$v3652\ := \$v3653\(4 to 35);
              case \$v3654\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11343_forever3163162\;
              when "0000" =>
                \$11351_i\ := \$v3652\(0 to 31);
                \$11338\ := \$11351_i\;
                \$v3651\ := \$$10700_pc_ptr_take\;
                if \$v3651\(0) = '1' then
                  state_var7021 <= q_wait3650;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr_write\ <= 0;
                  \$$10700_pc_write_request\ <= '1';
                  \$$10700_pc_write\ <= \$11338\;
                  state_var7021 <= pause_setI3648;
                end if;
              when others =>
                
              end case;
            when pause_getII3669 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11380\ := \$$10696_ram_value\;
              \$v3666\ := \$$10696_ram_ptr_take\;
              if \$v3666\(0) = '1' then
                state_var7021 <= q_wait3665;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11378_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11379\(0 to 35) & \$11331\(0 to 35) & \$11380\(72 to 107);
                state_var7021 <= pause_setI3663;
              end if;
            when pause_getII3676 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11379\ := \$$10696_ram_value\;
              \$v3672\ := "0000" & \$11330\;
              \$v3673\ := \$v3672\(0 to 3);
              \$v3667\ := \$v3672\(4 to 35);
              case \$v3673\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11398_forever3163165\;
              when "0000" =>
                \$11406_i\ := \$v3667\(0 to 31);
                \$v3671\ := \$$10696_ram_ptr_take\;
                if \$v3671\(0) = '1' then
                  state_var7021 <= q_wait3670;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11406_i\));
                  state_var7021 <= pause_getI3668;
                end if;
              when others =>
                
              end case;
            when pause_getII3685 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11331\ := \$$10696_ram_value\;
              \$v3681\ := "0000" & \$11330\;
              \$v3682\ := \$v3681\(0 to 3);
              \$v3662\ := \$v3681\(4 to 35);
              case \$v3682\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field1_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11370_forever3163164\;
              when "0000" =>
                \$11378_i\ := \$v3662\(0 to 31);
                \$v3679\ := "0000" & \$11330\;
                \$v3680\ := \$v3679\(0 to 3);
                \$v3674\ := \$v3679\(4 to 35);
                case \$v3680\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$11412_forever3163166\;
                when "0000" =>
                  \$11420_i\ := \$v3674\(0 to 31);
                  \$v3678\ := \$$10696_ram_ptr_take\;
                  if \$v3678\(0) = '1' then
                    state_var7021 <= q_wait3677;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$11420_i\));
                    state_var7021 <= pause_getI3675;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII3691 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11330\ := \$$10697_stack_value\;
              \$v3688\ := \$11328_cont\;
              \$v3689\ := \$v3688\(0 to 3);
              \$v3683\ := \$v3688\(4 to 35);
              case \$v3689\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11425_forever3163167\;
              when "0000" =>
                \$11433_i\ := \$v3683\(0 to 31);
                \$v3687\ := \$$10696_ram_ptr_take\;
                if \$v3687\(0) = '1' then
                  state_var7021 <= q_wait3686;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11433_i\));
                  state_var7021 <= pause_getI3684;
                end if;
              when others =>
                
              end case;
            when pause_getII3696 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11449\ := \$$10696_ram_value\;
              \$11437_loop3073170_arg\ := \$11449\(36 to 71) & eclat_unit;
              state_var7021 <= \$11437_loop3073170\;
            when pause_getII3707 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11443\ := \$$10696_ram_value\;
              \$v3703\ := \$11443\(72 to 107);
              \$v3704\ := \$v3703\(0 to 3);
              \$v3702\ := \$v3703\(4 to 35);
              case \$v3704\ is
              when "0001" =>
                \$11448\ := eclat_false;
              when "0000" =>
                \$11468_i\ := \$v3702\(0 to 31);
                \$11448\ := eclat_if(eclat_ge(\$11468_i\ & X"0000000" & X"0") & eclat_lt(\$11468_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3701\ := \$11448\;
              if \$v3701\(0) = '1' then
                \$11437_loop3073170_result\ := \$11437_loop3073170_arg\(0 to 35);
                \$11328_cont\ := \$11437_loop3073170_result\;
                \$v3693\ := \$$10697_stack_ptr_take\;
                if \$v3693\(0) = '1' then
                  state_var7021 <= q_wait3692;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3690;
                end if;
              else
                \$v3699\ := \$11437_loop3073170_arg\(0 to 35);
                \$v3700\ := \$v3699\(0 to 3);
                \$v3694\ := \$v3699\(4 to 35);
                case \$v3700\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$11458_forever3163168\;
                when "0000" =>
                  \$11466_i\ := \$v3694\(0 to 31);
                  \$v3698\ := \$$10696_ram_ptr_take\;
                  if \$v3698\(0) = '1' then
                    state_var7021 <= q_wait3697;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$11466_i\));
                    state_var7021 <= pause_getI3695;
                  end if;
                when others =>
                  
                end case;
              end if;
            when pause_getII3713 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11327\ := \$$10697_stack_value\;
              \$11437_loop3073170_arg\ := "0000" & \$11327\ & eclat_unit;
              state_var7021 <= \$11437_loop3073170\;
            when pause_getII3726 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11571\ := \$$10697_stack_value\;
              \$v3724\ := \$$10696_ram_ptr_take\;
              if \$v3724\(0) = '1' then
                state_var7021 <= q_wait3723;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3720\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11571\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11564_r\ & "0000" & \$11569\ & "0001" & \$v3720\;
                state_var7021 <= pause_setI3721;
              end if;
            when pause_getII3734 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11569\ := \$$10697_stack_value\;
              \$v3732\ := \$$10697_stack_ptr_take\;
              if \$v3732\(0) = '1' then
                state_var7021 <= q_wait3731;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11568_i\;
                state_var7021 <= pause_setI3729;
              end if;
            when pause_getII3738 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11568_i\ := \$$10702_brk_value\;
              \$v3736\ := \$$10697_stack_ptr_take\;
              if \$v3736\(0) = '1' then
                state_var7021 <= q_wait3735;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3733;
              end if;
            when pause_getII3742 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11568_i\ := \$$10702_brk_value\;
              \$v3736\ := \$$10697_stack_ptr_take\;
              if \$v3736\(0) = '1' then
                state_var7021 <= q_wait3735;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3733;
              end if;
            when pause_getII3750 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11576\ := \$$10702_brk_value\;
              \$v3748\ := \$$10702_brk_ptr_take\;
              if \$v3748\(0) = '1' then
                state_var7021 <= q_wait3747;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11576\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3745;
              end if;
            when pause_getII3755 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11567\ := \$$10695_limit_value\;
              \$v3753\ := eclat_eq(\$11566\ & eclat_sub(\$11567\ & X"0000000" & X"1"));
              if \$v3753\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11584_forever3163174\;
              else
                \$v3752\ := \$$10702_brk_ptr_take\;
                if \$v3752\(0) = '1' then
                  state_var7021 <= q_wait3751;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI3749;
                end if;
              end if;
            when pause_getII3759 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11566\ := \$$10702_brk_value\;
              \$v3757\ := \$$10695_limit_ptr_take\;
              if \$v3757\(0) = '1' then
                state_var7021 <= q_wait3756;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3754;
              end if;
            when pause_getII3763 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$11594\ := \$$10698_heap_value\;
              \$11564_r\ := "0000" & \$11594\;
              \$v3761\ := \$$10702_brk_ptr_take\;
              if \$v3761\(0) = '1' then
                state_var7021 <= q_wait3760;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3758;
              end if;
            when pause_getII3771 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$11562\ := \$$10698_heap_value\;
              \$v3769\ := \$$10696_ram_ptr_take\;
              if \$v3769\(0) = '1' then
                state_var7021 <= q_wait3768;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11562\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11556_z\ & \$11548_y\ & \$11540_x\;
                state_var7021 <= pause_setI3766;
              end if;
            when pause_getII3779 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11560_i\ := \$$10702_brk_value\;
              \$v3777\ := \$$10698_heap_ptr_take\;
              if \$v3777\(0) = '1' then
                state_var7021 <= q_wait3776;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11560_i\;
                state_var7021 <= pause_setI3774;
              end if;
            when pause_getII3783 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11560_i\ := \$$10702_brk_value\;
              \$v3777\ := \$$10698_heap_ptr_take\;
              if \$v3777\(0) = '1' then
                state_var7021 <= q_wait3776;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11560_i\;
                state_var7021 <= pause_setI3774;
              end if;
            when pause_getII3791 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11596\ := \$$10702_brk_value\;
              \$v3789\ := \$$10702_brk_ptr_take\;
              if \$v3789\(0) = '1' then
                state_var7021 <= q_wait3788;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11596\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3786;
              end if;
            when pause_getII3796 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11559\ := \$$10695_limit_value\;
              \$v3794\ := eclat_eq(\$11558\ & eclat_sub(\$11559\ & X"0000000" & X"1"));
              if \$v3794\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11604_forever3163175\;
              else
                \$v3793\ := \$$10702_brk_ptr_take\;
                if \$v3793\(0) = '1' then
                  state_var7021 <= q_wait3792;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI3790;
                end if;
              end if;
            when pause_getII3800 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11558\ := \$$10702_brk_value\;
              \$v3798\ := \$$10695_limit_ptr_take\;
              if \$v3798\(0) = '1' then
                state_var7021 <= q_wait3797;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3795;
              end if;
            when pause_getII3811 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11551\ := \$$10696_ram_value\;
              \$v3808\ := \$11551\(36 to 71);
              \$v3809\ := \$v3808\(0 to 3);
              \$v3807\ := \$v3808\(4 to 35);
              case \$v3809\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11619_forever3163176\;
              when "0000" =>
                \$11627_i\ := \$v3807\(0 to 31);
                \$11555\ := \$11627_i\;
                \$v3806\ := \$$10697_stack_ptr_take\;
                if \$v3806\(0) = '1' then
                  state_var7021 <= q_wait3805;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11555\;
                  state_var7021 <= pause_setI3803;
                end if;
              when others =>
                
              end case;
            when pause_getII3815 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11550\ := \$$10697_stack_value\;
              \$v3813\ := \$$10696_ram_ptr_take\;
              if \$v3813\(0) = '1' then
                state_var7021 <= q_wait3812;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11550\));
                state_var7021 <= pause_getI3810;
              end if;
            when pause_getII3826 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11543\ := \$$10696_ram_value\;
              \$v3823\ := \$11543\(36 to 71);
              \$v3824\ := \$v3823\(0 to 3);
              \$v3822\ := \$v3823\(4 to 35);
              case \$v3824\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11633_forever3163177\;
              when "0000" =>
                \$11641_i\ := \$v3822\(0 to 31);
                \$11547\ := \$11641_i\;
                \$v3821\ := \$$10697_stack_ptr_take\;
                if \$v3821\(0) = '1' then
                  state_var7021 <= q_wait3820;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11547\;
                  state_var7021 <= pause_setI3818;
                end if;
              when others =>
                
              end case;
            when pause_getII3830 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11542\ := \$$10697_stack_value\;
              \$v3828\ := \$$10696_ram_ptr_take\;
              if \$v3828\(0) = '1' then
                state_var7021 <= q_wait3827;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11542\));
                state_var7021 <= pause_getI3825;
              end if;
            when pause_getII3841 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11535\ := \$$10696_ram_value\;
              \$v3838\ := \$11535\(36 to 71);
              \$v3839\ := \$v3838\(0 to 3);
              \$v3837\ := \$v3838\(4 to 35);
              case \$v3839\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11647_forever3163178\;
              when "0000" =>
                \$11655_i\ := \$v3837\(0 to 31);
                \$11539\ := \$11655_i\;
                \$v3836\ := \$$10697_stack_ptr_take\;
                if \$v3836\(0) = '1' then
                  state_var7021 <= q_wait3835;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11539\;
                  state_var7021 <= pause_setI3833;
                end if;
              when others =>
                
              end case;
            when pause_getII3845 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11534\ := \$$10697_stack_value\;
              \$v3843\ := \$$10696_ram_ptr_take\;
              if \$v3843\(0) = '1' then
                state_var7021 <= q_wait3842;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11534\));
                state_var7021 <= pause_getI3840;
              end if;
            when pause_getII3854 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11670\ := \$$10697_stack_value\;
              \$v3852\ := \$$10696_ram_ptr_take\;
              if \$v3852\(0) = '1' then
                state_var7021 <= q_wait3851;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3848\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11670\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11663\ & "0000" & \$11668\ & "0001" & \$v3848\;
                state_var7021 <= pause_setI3849;
              end if;
            when pause_getII3862 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11668\ := \$$10697_stack_value\;
              \$v3860\ := \$$10697_stack_ptr_take\;
              if \$v3860\(0) = '1' then
                state_var7021 <= q_wait3859;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11667_i\;
                state_var7021 <= pause_setI3857;
              end if;
            when pause_getII3866 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11667_i\ := \$$10702_brk_value\;
              \$v3864\ := \$$10697_stack_ptr_take\;
              if \$v3864\(0) = '1' then
                state_var7021 <= q_wait3863;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3861;
              end if;
            when pause_getII3870 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11667_i\ := \$$10702_brk_value\;
              \$v3864\ := \$$10697_stack_ptr_take\;
              if \$v3864\(0) = '1' then
                state_var7021 <= q_wait3863;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3861;
              end if;
            when pause_getII3878 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11675\ := \$$10702_brk_value\;
              \$v3876\ := \$$10702_brk_ptr_take\;
              if \$v3876\(0) = '1' then
                state_var7021 <= q_wait3875;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11675\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3873;
              end if;
            when pause_getII3883 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11666\ := \$$10695_limit_value\;
              \$v3881\ := eclat_eq(\$11665\ & eclat_sub(\$11666\ & X"0000000" & X"1"));
              if \$v3881\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11683_forever3163179\;
              else
                \$v3880\ := \$$10702_brk_ptr_take\;
                if \$v3880\(0) = '1' then
                  state_var7021 <= q_wait3879;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI3877;
                end if;
              end if;
            when pause_getII3887 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11665\ := \$$10702_brk_value\;
              \$v3885\ := \$$10695_limit_ptr_take\;
              if \$v3885\(0) = '1' then
                state_var7021 <= q_wait3884;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3882;
              end if;
            when pause_getII3898 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11658\ := \$$10696_ram_value\;
              \$v3895\ := \$11658\(36 to 71);
              \$v3896\ := \$v3895\(0 to 3);
              \$v3894\ := \$v3895\(4 to 35);
              case \$v3896\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11698_forever3163180\;
              when "0000" =>
                \$11706_i\ := \$v3894\(0 to 31);
                \$11662\ := \$11706_i\;
                \$v3893\ := \$$10697_stack_ptr_take\;
                if \$v3893\(0) = '1' then
                  state_var7021 <= q_wait3892;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11662\;
                  state_var7021 <= pause_setI3890;
                end if;
              when others =>
                
              end case;
            when pause_getII3902 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11657\ := \$$10697_stack_value\;
              \$v3900\ := \$$10696_ram_ptr_take\;
              if \$v3900\(0) = '1' then
                state_var7021 <= q_wait3899;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11657\));
                state_var7021 <= pause_getI3897;
              end if;
            when pause_getII3913 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11709\ := \$$10696_ram_value\;
              \$v3910\ := \$11709\(36 to 71);
              \$v3911\ := \$v3910\(0 to 3);
              \$v3909\ := \$v3910\(4 to 35);
              case \$v3911\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11720_forever3163181\;
              when "0000" =>
                \$11728_i\ := \$v3909\(0 to 31);
                \$11713\ := \$11728_i\;
                \$v3908\ := \$$10697_stack_ptr_take\;
                if \$v3908\(0) = '1' then
                  state_var7021 <= q_wait3907;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11713\;
                  state_var7021 <= pause_setI3905;
                end if;
              when others =>
                
              end case;
            when pause_getII3917 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11708\ := \$$10697_stack_value\;
              \$v3915\ := \$$10696_ram_ptr_take\;
              if \$v3915\(0) = '1' then
                state_var7021 <= q_wait3914;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11708\));
                state_var7021 <= pause_getI3912;
              end if;
            when pause_getII3926 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11751\ := \$$10697_stack_value\;
              \$v3924\ := \$$10696_ram_ptr_take\;
              if \$v3924\(0) = '1' then
                state_var7021 <= q_wait3923;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3920\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11751\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11736_x\ & "0000" & \$11749\ & "0001" & \$v3920\;
                state_var7021 <= pause_setI3921;
              end if;
            when pause_getII3934 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11749\ := \$$10697_stack_value\;
              \$v3932\ := \$$10697_stack_ptr_take\;
              if \$v3932\(0) = '1' then
                state_var7021 <= q_wait3931;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11748_i\;
                state_var7021 <= pause_setI3929;
              end if;
            when pause_getII3938 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11748_i\ := \$$10702_brk_value\;
              \$v3936\ := \$$10697_stack_ptr_take\;
              if \$v3936\(0) = '1' then
                state_var7021 <= q_wait3935;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3933;
              end if;
            when pause_getII3942 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11748_i\ := \$$10702_brk_value\;
              \$v3936\ := \$$10697_stack_ptr_take\;
              if \$v3936\(0) = '1' then
                state_var7021 <= q_wait3935;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3933;
              end if;
            when pause_getII3950 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11756\ := \$$10702_brk_value\;
              \$v3948\ := \$$10702_brk_ptr_take\;
              if \$v3948\(0) = '1' then
                state_var7021 <= q_wait3947;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11756\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3945;
              end if;
            when pause_getII3955 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11747\ := \$$10695_limit_value\;
              \$v3953\ := eclat_eq(\$11746\ & eclat_sub(\$11747\ & X"0000000" & X"1"));
              if \$v3953\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11764_forever3163182\;
              else
                \$v3952\ := \$$10702_brk_ptr_take\;
                if \$v3952\(0) = '1' then
                  state_var7021 <= q_wait3951;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI3949;
                end if;
              end if;
            when pause_getII3959 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11746\ := \$$10702_brk_value\;
              \$v3957\ := \$$10695_limit_ptr_take\;
              if \$v3957\(0) = '1' then
                state_var7021 <= q_wait3956;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3954;
              end if;
            when pause_getII3970 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11739\ := \$$10696_ram_value\;
              \$v3967\ := \$11739\(36 to 71);
              \$v3968\ := \$v3967\(0 to 3);
              \$v3966\ := \$v3967\(4 to 35);
              case \$v3968\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11779_forever3163183\;
              when "0000" =>
                \$11787_i\ := \$v3966\(0 to 31);
                \$11743\ := \$11787_i\;
                \$v3965\ := \$$10697_stack_ptr_take\;
                if \$v3965\(0) = '1' then
                  state_var7021 <= q_wait3964;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11743\;
                  state_var7021 <= pause_setI3962;
                end if;
              when others =>
                
              end case;
            when pause_getII3974 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11738\ := \$$10697_stack_value\;
              \$v3972\ := \$$10696_ram_ptr_take\;
              if \$v3972\(0) = '1' then
                state_var7021 <= q_wait3971;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11738\));
                state_var7021 <= pause_getI3969;
              end if;
            when pause_getII3985 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11731\ := \$$10696_ram_value\;
              \$v3982\ := \$11731\(36 to 71);
              \$v3983\ := \$v3982\(0 to 3);
              \$v3981\ := \$v3982\(4 to 35);
              case \$v3983\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11793_forever3163184\;
              when "0000" =>
                \$11801_i\ := \$v3981\(0 to 31);
                \$11735\ := \$11801_i\;
                \$v3980\ := \$$10697_stack_ptr_take\;
                if \$v3980\(0) = '1' then
                  state_var7021 <= q_wait3979;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11735\;
                  state_var7021 <= pause_setI3977;
                end if;
              when others =>
                
              end case;
            when pause_getII3989 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11730\ := \$$10697_stack_value\;
              \$v3987\ := \$$10696_ram_ptr_take\;
              if \$v3987\(0) = '1' then
                state_var7021 <= q_wait3986;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11730\));
                state_var7021 <= pause_getI3984;
              end if;
            when pause_getII3998 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11821\ := \$$10697_stack_value\;
              \$v3996\ := \$$10696_ram_ptr_take\;
              if \$v3996\(0) = '1' then
                state_var7021 <= q_wait3995;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3992\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11821\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11814\ & "0000" & \$11819\ & "0001" & \$v3992\;
                state_var7021 <= pause_setI3993;
              end if;
            when pause_getII4006 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11819\ := \$$10697_stack_value\;
              \$v4004\ := \$$10697_stack_ptr_take\;
              if \$v4004\(0) = '1' then
                state_var7021 <= q_wait4003;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11818_i\;
                state_var7021 <= pause_setI4001;
              end if;
            when pause_getII4010 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11818_i\ := \$$10702_brk_value\;
              \$v4008\ := \$$10697_stack_ptr_take\;
              if \$v4008\(0) = '1' then
                state_var7021 <= q_wait4007;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4005;
              end if;
            when pause_getII4014 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11818_i\ := \$$10702_brk_value\;
              \$v4008\ := \$$10697_stack_ptr_take\;
              if \$v4008\(0) = '1' then
                state_var7021 <= q_wait4007;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4005;
              end if;
            when pause_getII4022 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11826\ := \$$10702_brk_value\;
              \$v4020\ := \$$10702_brk_ptr_take\;
              if \$v4020\(0) = '1' then
                state_var7021 <= q_wait4019;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11826\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4017;
              end if;
            when pause_getII4027 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11817\ := \$$10695_limit_value\;
              \$v4025\ := eclat_eq(\$11816\ & eclat_sub(\$11817\ & X"0000000" & X"1"));
              if \$v4025\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11834_forever3163185\;
              else
                \$v4024\ := \$$10702_brk_ptr_take\;
                if \$v4024\(0) = '1' then
                  state_var7021 <= q_wait4023;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4021;
                end if;
              end if;
            when pause_getII4031 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11816\ := \$$10702_brk_value\;
              \$v4029\ := \$$10695_limit_ptr_take\;
              if \$v4029\(0) = '1' then
                state_var7021 <= q_wait4028;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4026;
              end if;
            when pause_getII4035 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$11854\ := \$$10698_heap_value\;
              \$11814\ := "0000" & \$11854\;
              \$v4033\ := \$$10702_brk_ptr_take\;
              if \$v4033\(0) = '1' then
                state_var7021 <= q_wait4032;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4030;
              end if;
            when pause_getII4044 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$11848\ := \$$10698_heap_value\;
              \$v4042\ := \$$10696_ram_ptr_take\;
              if \$v4042\(0) = '1' then
                state_var7021 <= q_wait4041;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4038\ := X"0000000" & X"1";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11848\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11810\(0 to 35) & "0000" & \$11812\ & "0001" & \$v4038\;
                state_var7021 <= pause_setI4039;
              end if;
            when pause_getII4052 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11846_i\ := \$$10702_brk_value\;
              \$v4050\ := \$$10698_heap_ptr_take\;
              if \$v4050\(0) = '1' then
                state_var7021 <= q_wait4049;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11846_i\;
                state_var7021 <= pause_setI4047;
              end if;
            when pause_getII4056 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11846_i\ := \$$10702_brk_value\;
              \$v4050\ := \$$10698_heap_ptr_take\;
              if \$v4050\(0) = '1' then
                state_var7021 <= q_wait4049;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11846_i\;
                state_var7021 <= pause_setI4047;
              end if;
            when pause_getII4064 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11859\ := \$$10702_brk_value\;
              \$v4062\ := \$$10702_brk_ptr_take\;
              if \$v4062\(0) = '1' then
                state_var7021 <= q_wait4061;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11859\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4059;
              end if;
            when pause_getII4069 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11845\ := \$$10695_limit_value\;
              \$v4067\ := eclat_eq(\$11844\ & eclat_sub(\$11845\ & X"0000000" & X"1"));
              if \$v4067\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11867_forever3163186\;
              else
                \$v4066\ := \$$10702_brk_ptr_take\;
                if \$v4066\(0) = '1' then
                  state_var7021 <= q_wait4065;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4063;
                end if;
              end if;
            when pause_getII4073 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11844\ := \$$10702_brk_value\;
              \$v4071\ := \$$10695_limit_ptr_take\;
              if \$v4071\(0) = '1' then
                state_var7021 <= q_wait4070;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4068;
              end if;
            when pause_getII4077 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11812\ := \$$10697_stack_value\;
              \$v4075\ := \$$10702_brk_ptr_take\;
              if \$v4075\(0) = '1' then
                state_var7021 <= q_wait4074;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4072;
              end if;
            when pause_getII4082 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11810\ := \$$10696_ram_value\;
              \$v4079\ := \$$10697_stack_ptr_take\;
              if \$v4079\(0) = '1' then
                state_var7021 <= q_wait4078;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4076;
              end if;
            when pause_getII4095 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11804\ := \$$10696_ram_value\;
              \$v4092\ := \$11804\(36 to 71);
              \$v4093\ := \$v4092\(0 to 3);
              \$v4091\ := \$v4092\(4 to 35);
              case \$v4093\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11895_forever3163188\;
              when "0000" =>
                \$11903_i\ := \$v4091\(0 to 31);
                \$11808\ := \$11903_i\;
                \$v4090\ := \$$10697_stack_ptr_take\;
                if \$v4090\(0) = '1' then
                  state_var7021 <= q_wait4089;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11808\;
                  state_var7021 <= pause_setI4087;
                end if;
              when others =>
                
              end case;
            when pause_getII4099 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11803\ := \$$10697_stack_value\;
              \$v4097\ := \$$10696_ram_ptr_take\;
              if \$v4097\(0) = '1' then
                state_var7021 <= q_wait4096;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11803\));
                state_var7021 <= pause_getI4094;
              end if;
            when pause_getII4110 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11919\ := \$$10697_stack_value\;
              \$v4108\ := \$$10696_ram_ptr_take\;
              if \$v4108\(0) = '1' then
                state_var7021 <= q_wait4107;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4103\ := X"0000000" & X"1";
                \$v4102\ := X"0000000" & X"2";
                \$v4104\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11919\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= eclat_if(\$11912\ & "0000" & \$v4103\ & "0000" & \$v4102\) & "0000" & \$11917\ & "0001" & \$v4104\;
                state_var7021 <= pause_setI4105;
              end if;
            when pause_getII4118 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11917\ := \$$10697_stack_value\;
              \$v4116\ := \$$10697_stack_ptr_take\;
              if \$v4116\(0) = '1' then
                state_var7021 <= q_wait4115;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11916_i\;
                state_var7021 <= pause_setI4113;
              end if;
            when pause_getII4122 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11916_i\ := \$$10702_brk_value\;
              \$v4120\ := \$$10697_stack_ptr_take\;
              if \$v4120\(0) = '1' then
                state_var7021 <= q_wait4119;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4117;
              end if;
            when pause_getII4126 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11916_i\ := \$$10702_brk_value\;
              \$v4120\ := \$$10697_stack_ptr_take\;
              if \$v4120\(0) = '1' then
                state_var7021 <= q_wait4119;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4117;
              end if;
            when pause_getII4134 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11925\ := \$$10702_brk_value\;
              \$v4132\ := \$$10702_brk_ptr_take\;
              if \$v4132\(0) = '1' then
                state_var7021 <= q_wait4131;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11925\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4129;
              end if;
            when pause_getII4139 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11915\ := \$$10695_limit_value\;
              \$v4137\ := eclat_eq(\$11914\ & eclat_sub(\$11915\ & X"0000000" & X"1"));
              if \$v4137\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11933_forever3163189\;
              else
                \$v4136\ := \$$10702_brk_ptr_take\;
                if \$v4136\(0) = '1' then
                  state_var7021 <= q_wait4135;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4133;
                end if;
              end if;
            when pause_getII4143 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11914\ := \$$10702_brk_value\;
              \$v4141\ := \$$10695_limit_ptr_take\;
              if \$v4141\(0) = '1' then
                state_var7021 <= q_wait4140;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4138;
              end if;
            when pause_getII4157 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11906\ := \$$10696_ram_value\;
              \$v4154\ := \$11906\(36 to 71);
              \$v4155\ := \$v4154\(0 to 3);
              \$v4153\ := \$v4154\(4 to 35);
              case \$v4155\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11951_forever3163190\;
              when "0000" =>
                \$11959_i\ := \$v4153\(0 to 31);
                \$11910\ := \$11959_i\;
                \$v4152\ := \$$10697_stack_ptr_take\;
                if \$v4152\(0) = '1' then
                  state_var7021 <= q_wait4151;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11910\;
                  state_var7021 <= pause_setI4149;
                end if;
              when others =>
                
              end case;
            when pause_getII4161 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11905\ := \$$10697_stack_value\;
              \$v4159\ := \$$10696_ram_ptr_take\;
              if \$v4159\(0) = '1' then
                state_var7021 <= q_wait4158;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11905\));
                state_var7021 <= pause_getI4156;
              end if;
            when pause_getII4170 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11975\ := \$$10697_stack_value\;
              \$v4168\ := \$$10696_ram_ptr_take\;
              if \$v4168\(0) = '1' then
                state_var7021 <= q_wait4167;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4164\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11975\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11968\(0 to 35) & "0000" & \$11973\ & "0001" & \$v4164\;
                state_var7021 <= pause_setI4165;
              end if;
            when pause_getII4178 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11973\ := \$$10697_stack_value\;
              \$v4176\ := \$$10697_stack_ptr_take\;
              if \$v4176\(0) = '1' then
                state_var7021 <= q_wait4175;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11972_i\;
                state_var7021 <= pause_setI4173;
              end if;
            when pause_getII4182 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11972_i\ := \$$10702_brk_value\;
              \$v4180\ := \$$10697_stack_ptr_take\;
              if \$v4180\(0) = '1' then
                state_var7021 <= q_wait4179;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4177;
              end if;
            when pause_getII4186 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11972_i\ := \$$10702_brk_value\;
              \$v4180\ := \$$10697_stack_ptr_take\;
              if \$v4180\(0) = '1' then
                state_var7021 <= q_wait4179;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4177;
              end if;
            when pause_getII4194 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11984\ := \$$10702_brk_value\;
              \$v4192\ := \$$10702_brk_ptr_take\;
              if \$v4192\(0) = '1' then
                state_var7021 <= q_wait4191;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11984\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4189;
              end if;
            when pause_getII4199 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$11971\ := \$$10695_limit_value\;
              \$v4197\ := eclat_eq(\$11970\ & eclat_sub(\$11971\ & X"0000000" & X"1"));
              if \$v4197\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11992_forever3163191\;
              else
                \$v4196\ := \$$10702_brk_ptr_take\;
                if \$v4196\(0) = '1' then
                  state_var7021 <= q_wait4195;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4193;
                end if;
              end if;
            when pause_getII4203 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$11970\ := \$$10702_brk_value\;
              \$v4201\ := \$$10695_limit_ptr_take\;
              if \$v4201\(0) = '1' then
                state_var7021 <= q_wait4200;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4198;
              end if;
            when pause_getII4208 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11968\ := \$$10696_ram_value\;
              \$v4205\ := \$$10702_brk_ptr_take\;
              if \$v4205\(0) = '1' then
                state_var7021 <= q_wait4204;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4202;
              end if;
            when pause_getII4221 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$11962\ := \$$10696_ram_value\;
              \$v4218\ := \$11962\(36 to 71);
              \$v4219\ := \$v4218\(0 to 3);
              \$v4217\ := \$v4218\(4 to 35);
              case \$v4219\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12020_forever3163193\;
              when "0000" =>
                \$12028_i\ := \$v4217\(0 to 31);
                \$11966\ := \$12028_i\;
                \$v4216\ := \$$10697_stack_ptr_take\;
                if \$v4216\(0) = '1' then
                  state_var7021 <= q_wait4215;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$11966\;
                  state_var7021 <= pause_setI4213;
                end if;
              when others =>
                
              end case;
            when pause_getII4225 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11961\ := \$$10697_stack_value\;
              \$v4223\ := \$$10696_ram_ptr_take\;
              if \$v4223\(0) = '1' then
                state_var7021 <= q_wait4222;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11961\));
                state_var7021 <= pause_getI4220;
              end if;
            when pause_getII4234 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12044\ := \$$10697_stack_value\;
              \$v4232\ := \$$10696_ram_ptr_take\;
              if \$v4232\(0) = '1' then
                state_var7021 <= q_wait4231;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4228\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12044\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12037\(36 to 71) & "0000" & \$12042\ & "0001" & \$v4228\;
                state_var7021 <= pause_setI4229;
              end if;
            when pause_getII4242 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12042\ := \$$10697_stack_value\;
              \$v4240\ := \$$10697_stack_ptr_take\;
              if \$v4240\(0) = '1' then
                state_var7021 <= q_wait4239;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12041_i\;
                state_var7021 <= pause_setI4237;
              end if;
            when pause_getII4246 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12041_i\ := \$$10702_brk_value\;
              \$v4244\ := \$$10697_stack_ptr_take\;
              if \$v4244\(0) = '1' then
                state_var7021 <= q_wait4243;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4241;
              end if;
            when pause_getII4250 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12041_i\ := \$$10702_brk_value\;
              \$v4244\ := \$$10697_stack_ptr_take\;
              if \$v4244\(0) = '1' then
                state_var7021 <= q_wait4243;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4241;
              end if;
            when pause_getII4258 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12053\ := \$$10702_brk_value\;
              \$v4256\ := \$$10702_brk_ptr_take\;
              if \$v4256\(0) = '1' then
                state_var7021 <= q_wait4255;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12053\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4253;
              end if;
            when pause_getII4263 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12040\ := \$$10695_limit_value\;
              \$v4261\ := eclat_eq(\$12039\ & eclat_sub(\$12040\ & X"0000000" & X"1"));
              if \$v4261\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12061_forever3163194\;
              else
                \$v4260\ := \$$10702_brk_ptr_take\;
                if \$v4260\(0) = '1' then
                  state_var7021 <= q_wait4259;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4257;
                end if;
              end if;
            when pause_getII4267 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12039\ := \$$10702_brk_value\;
              \$v4265\ := \$$10695_limit_ptr_take\;
              if \$v4265\(0) = '1' then
                state_var7021 <= q_wait4264;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4262;
              end if;
            when pause_getII4272 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12037\ := \$$10696_ram_value\;
              \$v4269\ := \$$10702_brk_ptr_take\;
              if \$v4269\(0) = '1' then
                state_var7021 <= q_wait4268;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4266;
              end if;
            when pause_getII4285 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12031\ := \$$10696_ram_value\;
              \$v4282\ := \$12031\(36 to 71);
              \$v4283\ := \$v4282\(0 to 3);
              \$v4281\ := \$v4282\(4 to 35);
              case \$v4283\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12089_forever3163196\;
              when "0000" =>
                \$12097_i\ := \$v4281\(0 to 31);
                \$12035\ := \$12097_i\;
                \$v4280\ := \$$10697_stack_ptr_take\;
                if \$v4280\(0) = '1' then
                  state_var7021 <= q_wait4279;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12035\;
                  state_var7021 <= pause_setI4277;
                end if;
              when others =>
                
              end case;
            when pause_getII4289 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12030\ := \$$10697_stack_value\;
              \$v4287\ := \$$10696_ram_ptr_take\;
              if \$v4287\(0) = '1' then
                state_var7021 <= q_wait4286;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12030\));
                state_var7021 <= pause_getI4284;
              end if;
            when pause_getII4298 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12113\ := \$$10697_stack_value\;
              \$v4296\ := \$$10696_ram_ptr_take\;
              if \$v4296\(0) = '1' then
                state_var7021 <= q_wait4295;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4292\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12113\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12106\(72 to 107) & "0000" & \$12111\ & "0001" & \$v4292\;
                state_var7021 <= pause_setI4293;
              end if;
            when pause_getII4306 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12111\ := \$$10697_stack_value\;
              \$v4304\ := \$$10697_stack_ptr_take\;
              if \$v4304\(0) = '1' then
                state_var7021 <= q_wait4303;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12110_i\;
                state_var7021 <= pause_setI4301;
              end if;
            when pause_getII4310 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12110_i\ := \$$10702_brk_value\;
              \$v4308\ := \$$10697_stack_ptr_take\;
              if \$v4308\(0) = '1' then
                state_var7021 <= q_wait4307;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4305;
              end if;
            when pause_getII4314 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12110_i\ := \$$10702_brk_value\;
              \$v4308\ := \$$10697_stack_ptr_take\;
              if \$v4308\(0) = '1' then
                state_var7021 <= q_wait4307;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4305;
              end if;
            when pause_getII4322 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12122\ := \$$10702_brk_value\;
              \$v4320\ := \$$10702_brk_ptr_take\;
              if \$v4320\(0) = '1' then
                state_var7021 <= q_wait4319;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12122\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4317;
              end if;
            when pause_getII4327 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12109\ := \$$10695_limit_value\;
              \$v4325\ := eclat_eq(\$12108\ & eclat_sub(\$12109\ & X"0000000" & X"1"));
              if \$v4325\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12130_forever3163197\;
              else
                \$v4324\ := \$$10702_brk_ptr_take\;
                if \$v4324\(0) = '1' then
                  state_var7021 <= q_wait4323;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4321;
                end if;
              end if;
            when pause_getII4331 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12108\ := \$$10702_brk_value\;
              \$v4329\ := \$$10695_limit_ptr_take\;
              if \$v4329\(0) = '1' then
                state_var7021 <= q_wait4328;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4326;
              end if;
            when pause_getII4336 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12106\ := \$$10696_ram_value\;
              \$v4333\ := \$$10702_brk_ptr_take\;
              if \$v4333\(0) = '1' then
                state_var7021 <= q_wait4332;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4330;
              end if;
            when pause_getII4349 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12100\ := \$$10696_ram_value\;
              \$v4346\ := \$12100\(36 to 71);
              \$v4347\ := \$v4346\(0 to 3);
              \$v4345\ := \$v4346\(4 to 35);
              case \$v4347\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12158_forever3163199\;
              when "0000" =>
                \$12166_i\ := \$v4345\(0 to 31);
                \$12104\ := \$12166_i\;
                \$v4344\ := \$$10697_stack_ptr_take\;
                if \$v4344\(0) = '1' then
                  state_var7021 <= q_wait4343;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12104\;
                  state_var7021 <= pause_setI4341;
                end if;
              when others =>
                
              end case;
            when pause_getII4353 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12099\ := \$$10697_stack_value\;
              \$v4351\ := \$$10696_ram_ptr_take\;
              if \$v4351\(0) = '1' then
                state_var7021 <= q_wait4350;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12099\));
                state_var7021 <= pause_getI4348;
              end if;
            when pause_getII4362 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12190\ := \$$10697_stack_value\;
              \$v4360\ := \$$10696_ram_ptr_take\;
              if \$v4360\(0) = '1' then
                state_var7021 <= q_wait4359;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4356\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12190\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12174_x\ & "0000" & \$12188\ & "0001" & \$v4356\;
                state_var7021 <= pause_setI4357;
              end if;
            when pause_getII4370 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12188\ := \$$10697_stack_value\;
              \$v4368\ := \$$10697_stack_ptr_take\;
              if \$v4368\(0) = '1' then
                state_var7021 <= q_wait4367;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12187_i\;
                state_var7021 <= pause_setI4365;
              end if;
            when pause_getII4374 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12187_i\ := \$$10702_brk_value\;
              \$v4372\ := \$$10697_stack_ptr_take\;
              if \$v4372\(0) = '1' then
                state_var7021 <= q_wait4371;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4369;
              end if;
            when pause_getII4378 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12187_i\ := \$$10702_brk_value\;
              \$v4372\ := \$$10697_stack_ptr_take\;
              if \$v4372\(0) = '1' then
                state_var7021 <= q_wait4371;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4369;
              end if;
            when pause_getII4386 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12195\ := \$$10702_brk_value\;
              \$v4384\ := \$$10702_brk_ptr_take\;
              if \$v4384\(0) = '1' then
                state_var7021 <= q_wait4383;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12195\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4381;
              end if;
            when pause_getII4391 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12186\ := \$$10695_limit_value\;
              \$v4389\ := eclat_eq(\$12185\ & eclat_sub(\$12186\ & X"0000000" & X"1"));
              if \$v4389\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12203_forever3163200\;
              else
                \$v4388\ := \$$10702_brk_ptr_take\;
                if \$v4388\(0) = '1' then
                  state_var7021 <= q_wait4387;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4385;
                end if;
              end if;
            when pause_getII4395 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12185\ := \$$10702_brk_value\;
              \$v4393\ := \$$10695_limit_ptr_take\;
              if \$v4393\(0) = '1' then
                state_var7021 <= q_wait4392;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4390;
              end if;
            when pause_getII4405 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12227\ := \$$10696_ram_value\;
              \$v4402\ := \$$10696_ram_ptr_take\;
              if \$v4402\(0) = '1' then
                state_var7021 <= q_wait4401;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12225_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12174_x\ & \$12226\(36 to 71) & \$12227\(72 to 107);
                state_var7021 <= pause_setI4399;
              end if;
            when pause_getII4412 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12226\ := \$$10696_ram_value\;
              \$v4408\ := \$12182_y\;
              \$v4409\ := \$v4408\(0 to 3);
              \$v4403\ := \$v4408\(4 to 35);
              case \$v4409\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12240_forever3163202\;
              when "0000" =>
                \$12248_i\ := \$v4403\(0 to 31);
                \$v4407\ := \$$10696_ram_ptr_take\;
                if \$v4407\(0) = '1' then
                  state_var7021 <= q_wait4406;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$12248_i\));
                  state_var7021 <= pause_getI4404;
                end if;
              when others =>
                
              end case;
            when pause_getII4427 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12177\ := \$$10696_ram_value\;
              \$v4424\ := \$12177\(36 to 71);
              \$v4425\ := \$v4424\(0 to 3);
              \$v4423\ := \$v4424\(4 to 35);
              case \$v4425\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12267_forever3163204\;
              when "0000" =>
                \$12275_i\ := \$v4423\(0 to 31);
                \$12181\ := \$12275_i\;
                \$v4422\ := \$$10697_stack_ptr_take\;
                if \$v4422\(0) = '1' then
                  state_var7021 <= q_wait4421;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12181\;
                  state_var7021 <= pause_setI4419;
                end if;
              when others =>
                
              end case;
            when pause_getII4431 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12176\ := \$$10697_stack_value\;
              \$v4429\ := \$$10696_ram_ptr_take\;
              if \$v4429\(0) = '1' then
                state_var7021 <= q_wait4428;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12176\));
                state_var7021 <= pause_getI4426;
              end if;
            when pause_getII4442 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12169\ := \$$10696_ram_value\;
              \$v4439\ := \$12169\(36 to 71);
              \$v4440\ := \$v4439\(0 to 3);
              \$v4438\ := \$v4439\(4 to 35);
              case \$v4440\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12281_forever3163205\;
              when "0000" =>
                \$12289_i\ := \$v4438\(0 to 31);
                \$12173\ := \$12289_i\;
                \$v4437\ := \$$10697_stack_ptr_take\;
                if \$v4437\(0) = '1' then
                  state_var7021 <= q_wait4436;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12173\;
                  state_var7021 <= pause_setI4434;
                end if;
              when others =>
                
              end case;
            when pause_getII4446 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12168\ := \$$10697_stack_value\;
              \$v4444\ := \$$10696_ram_ptr_take\;
              if \$v4444\(0) = '1' then
                state_var7021 <= q_wait4443;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12168\));
                state_var7021 <= pause_getI4441;
              end if;
            when pause_getII4455 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12313\ := \$$10697_stack_value\;
              \$v4453\ := \$$10696_ram_ptr_take\;
              if \$v4453\(0) = '1' then
                state_var7021 <= q_wait4452;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4449\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12313\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12297_x\ & "0000" & \$12311\ & "0001" & \$v4449\;
                state_var7021 <= pause_setI4450;
              end if;
            when pause_getII4463 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12311\ := \$$10697_stack_value\;
              \$v4461\ := \$$10697_stack_ptr_take\;
              if \$v4461\(0) = '1' then
                state_var7021 <= q_wait4460;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12310_i\;
                state_var7021 <= pause_setI4458;
              end if;
            when pause_getII4467 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12310_i\ := \$$10702_brk_value\;
              \$v4465\ := \$$10697_stack_ptr_take\;
              if \$v4465\(0) = '1' then
                state_var7021 <= q_wait4464;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4462;
              end if;
            when pause_getII4471 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12310_i\ := \$$10702_brk_value\;
              \$v4465\ := \$$10697_stack_ptr_take\;
              if \$v4465\(0) = '1' then
                state_var7021 <= q_wait4464;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4462;
              end if;
            when pause_getII4479 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12318\ := \$$10702_brk_value\;
              \$v4477\ := \$$10702_brk_ptr_take\;
              if \$v4477\(0) = '1' then
                state_var7021 <= q_wait4476;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12318\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4474;
              end if;
            when pause_getII4484 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12309\ := \$$10695_limit_value\;
              \$v4482\ := eclat_eq(\$12308\ & eclat_sub(\$12309\ & X"0000000" & X"1"));
              if \$v4482\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12326_forever3163206\;
              else
                \$v4481\ := \$$10702_brk_ptr_take\;
                if \$v4481\(0) = '1' then
                  state_var7021 <= q_wait4480;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4478;
                end if;
              end if;
            when pause_getII4488 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12308\ := \$$10702_brk_value\;
              \$v4486\ := \$$10695_limit_ptr_take\;
              if \$v4486\(0) = '1' then
                state_var7021 <= q_wait4485;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4483;
              end if;
            when pause_getII4498 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12350\ := \$$10696_ram_value\;
              \$v4495\ := \$$10696_ram_ptr_take\;
              if \$v4495\(0) = '1' then
                state_var7021 <= q_wait4494;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12348_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12349\(0 to 35) & \$12297_x\ & \$12350\(72 to 107);
                state_var7021 <= pause_setI4492;
              end if;
            when pause_getII4505 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12349\ := \$$10696_ram_value\;
              \$v4501\ := \$12305_y\;
              \$v4502\ := \$v4501\(0 to 3);
              \$v4496\ := \$v4501\(4 to 35);
              case \$v4502\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12363_forever3163208\;
              when "0000" =>
                \$12371_i\ := \$v4496\(0 to 31);
                \$v4500\ := \$$10696_ram_ptr_take\;
                if \$v4500\(0) = '1' then
                  state_var7021 <= q_wait4499;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$12371_i\));
                  state_var7021 <= pause_getI4497;
                end if;
              when others =>
                
              end case;
            when pause_getII4520 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12300\ := \$$10696_ram_value\;
              \$v4517\ := \$12300\(36 to 71);
              \$v4518\ := \$v4517\(0 to 3);
              \$v4516\ := \$v4517\(4 to 35);
              case \$v4518\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12390_forever3163210\;
              when "0000" =>
                \$12398_i\ := \$v4516\(0 to 31);
                \$12304\ := \$12398_i\;
                \$v4515\ := \$$10697_stack_ptr_take\;
                if \$v4515\(0) = '1' then
                  state_var7021 <= q_wait4514;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12304\;
                  state_var7021 <= pause_setI4512;
                end if;
              when others =>
                
              end case;
            when pause_getII4524 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12299\ := \$$10697_stack_value\;
              \$v4522\ := \$$10696_ram_ptr_take\;
              if \$v4522\(0) = '1' then
                state_var7021 <= q_wait4521;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12299\));
                state_var7021 <= pause_getI4519;
              end if;
            when pause_getII4535 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12292\ := \$$10696_ram_value\;
              \$v4532\ := \$12292\(36 to 71);
              \$v4533\ := \$v4532\(0 to 3);
              \$v4531\ := \$v4532\(4 to 35);
              case \$v4533\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12404_forever3163211\;
              when "0000" =>
                \$12412_i\ := \$v4531\(0 to 31);
                \$12296\ := \$12412_i\;
                \$v4530\ := \$$10697_stack_ptr_take\;
                if \$v4530\(0) = '1' then
                  state_var7021 <= q_wait4529;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12296\;
                  state_var7021 <= pause_setI4527;
                end if;
              when others =>
                
              end case;
            when pause_getII4539 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12291\ := \$$10697_stack_value\;
              \$v4537\ := \$$10696_ram_ptr_take\;
              if \$v4537\(0) = '1' then
                state_var7021 <= q_wait4536;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12291\));
                state_var7021 <= pause_getI4534;
              end if;
            when pause_getII4548 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12436\ := \$$10697_stack_value\;
              \$v4546\ := \$$10696_ram_ptr_take\;
              if \$v4546\(0) = '1' then
                state_var7021 <= q_wait4545;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4542\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12436\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12420_x\ & "0000" & \$12434\ & "0001" & \$v4542\;
                state_var7021 <= pause_setI4543;
              end if;
            when pause_getII4556 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12434\ := \$$10697_stack_value\;
              \$v4554\ := \$$10697_stack_ptr_take\;
              if \$v4554\(0) = '1' then
                state_var7021 <= q_wait4553;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12433_i\;
                state_var7021 <= pause_setI4551;
              end if;
            when pause_getII4560 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12433_i\ := \$$10702_brk_value\;
              \$v4558\ := \$$10697_stack_ptr_take\;
              if \$v4558\(0) = '1' then
                state_var7021 <= q_wait4557;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4555;
              end if;
            when pause_getII4564 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12433_i\ := \$$10702_brk_value\;
              \$v4558\ := \$$10697_stack_ptr_take\;
              if \$v4558\(0) = '1' then
                state_var7021 <= q_wait4557;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4555;
              end if;
            when pause_getII4572 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12441\ := \$$10702_brk_value\;
              \$v4570\ := \$$10702_brk_ptr_take\;
              if \$v4570\(0) = '1' then
                state_var7021 <= q_wait4569;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12441\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4567;
              end if;
            when pause_getII4577 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12432\ := \$$10695_limit_value\;
              \$v4575\ := eclat_eq(\$12431\ & eclat_sub(\$12432\ & X"0000000" & X"1"));
              if \$v4575\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12449_forever3163212\;
              else
                \$v4574\ := \$$10702_brk_ptr_take\;
                if \$v4574\(0) = '1' then
                  state_var7021 <= q_wait4573;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4571;
                end if;
              end if;
            when pause_getII4581 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12431\ := \$$10702_brk_value\;
              \$v4579\ := \$$10695_limit_ptr_take\;
              if \$v4579\(0) = '1' then
                state_var7021 <= q_wait4578;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4576;
              end if;
            when pause_getII4591 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12473\ := \$$10696_ram_value\;
              \$v4588\ := \$$10696_ram_ptr_take\;
              if \$v4588\(0) = '1' then
                state_var7021 <= q_wait4587;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12471_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12472\(0 to 35) & \$12473\(36 to 71) & \$12420_x\;
                state_var7021 <= pause_setI4585;
              end if;
            when pause_getII4598 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12472\ := \$$10696_ram_value\;
              \$v4594\ := \$12428_y\;
              \$v4595\ := \$v4594\(0 to 3);
              \$v4589\ := \$v4594\(4 to 35);
              case \$v4595\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12486_forever3163214\;
              when "0000" =>
                \$12494_i\ := \$v4589\(0 to 31);
                \$v4593\ := \$$10696_ram_ptr_take\;
                if \$v4593\(0) = '1' then
                  state_var7021 <= q_wait4592;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$12494_i\));
                  state_var7021 <= pause_getI4590;
                end if;
              when others =>
                
              end case;
            when pause_getII4613 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12423\ := \$$10696_ram_value\;
              \$v4610\ := \$12423\(36 to 71);
              \$v4611\ := \$v4610\(0 to 3);
              \$v4609\ := \$v4610\(4 to 35);
              case \$v4611\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12513_forever3163216\;
              when "0000" =>
                \$12521_i\ := \$v4609\(0 to 31);
                \$12427\ := \$12521_i\;
                \$v4608\ := \$$10697_stack_ptr_take\;
                if \$v4608\(0) = '1' then
                  state_var7021 <= q_wait4607;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12427\;
                  state_var7021 <= pause_setI4605;
                end if;
              when others =>
                
              end case;
            when pause_getII4617 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12422\ := \$$10697_stack_value\;
              \$v4615\ := \$$10696_ram_ptr_take\;
              if \$v4615\(0) = '1' then
                state_var7021 <= q_wait4614;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12422\));
                state_var7021 <= pause_getI4612;
              end if;
            when pause_getII4628 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12415\ := \$$10696_ram_value\;
              \$v4625\ := \$12415\(36 to 71);
              \$v4626\ := \$v4625\(0 to 3);
              \$v4624\ := \$v4625\(4 to 35);
              case \$v4626\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12527_forever3163217\;
              when "0000" =>
                \$12535_i\ := \$v4624\(0 to 31);
                \$12419\ := \$12535_i\;
                \$v4623\ := \$$10697_stack_ptr_take\;
                if \$v4623\(0) = '1' then
                  state_var7021 <= q_wait4622;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12419\;
                  state_var7021 <= pause_setI4620;
                end if;
              when others =>
                
              end case;
            when pause_getII4632 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12414\ := \$$10697_stack_value\;
              \$v4630\ := \$$10696_ram_ptr_take\;
              if \$v4630\(0) = '1' then
                state_var7021 <= q_wait4629;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12414\));
                state_var7021 <= pause_getI4627;
              end if;
            when pause_getII4643 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12559\ := \$$10697_stack_value\;
              \$v4641\ := \$$10696_ram_ptr_take\;
              if \$v4641\(0) = '1' then
                state_var7021 <= q_wait4640;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4636\ := X"0000000" & X"1";
                \$v4635\ := X"0000000" & X"2";
                \$v4637\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12559\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= eclat_if(\$12552\ & "0000" & \$v4636\ & "0000" & \$v4635\) & "0000" & \$12557\ & "0001" & \$v4637\;
                state_var7021 <= pause_setI4638;
              end if;
            when pause_getII4651 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12557\ := \$$10697_stack_value\;
              \$v4649\ := \$$10697_stack_ptr_take\;
              if \$v4649\(0) = '1' then
                state_var7021 <= q_wait4648;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12556_i\;
                state_var7021 <= pause_setI4646;
              end if;
            when pause_getII4655 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12556_i\ := \$$10702_brk_value\;
              \$v4653\ := \$$10697_stack_ptr_take\;
              if \$v4653\(0) = '1' then
                state_var7021 <= q_wait4652;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4650;
              end if;
            when pause_getII4659 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12556_i\ := \$$10702_brk_value\;
              \$v4653\ := \$$10697_stack_ptr_take\;
              if \$v4653\(0) = '1' then
                state_var7021 <= q_wait4652;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4650;
              end if;
            when pause_getII4667 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12565\ := \$$10702_brk_value\;
              \$v4665\ := \$$10702_brk_ptr_take\;
              if \$v4665\(0) = '1' then
                state_var7021 <= q_wait4664;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12565\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4662;
              end if;
            when pause_getII4672 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12555\ := \$$10695_limit_value\;
              \$v4670\ := eclat_eq(\$12554\ & eclat_sub(\$12555\ & X"0000000" & X"1"));
              if \$v4670\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12573_forever3163218\;
              else
                \$v4669\ := \$$10702_brk_ptr_take\;
                if \$v4669\(0) = '1' then
                  state_var7021 <= q_wait4668;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4666;
                end if;
              end if;
            when pause_getII4676 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12554\ := \$$10702_brk_value\;
              \$v4674\ := \$$10695_limit_ptr_take\;
              if \$v4674\(0) = '1' then
                state_var7021 <= q_wait4673;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4671;
              end if;
            when pause_getII4715 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12588\ := \$$10696_ram_value\;
              \$v4711\ := \$12587\(0 to 35);
              \$v4712\ := \$v4711\(0 to 3);
              \$v4704\ := \$v4711\(4 to 35);
              case \$v4712\ is
              when "0001" =>
                \$12611_i\ := \$v4704\(0 to 31);
                \$v4706\ := \$12588\(0 to 35);
                \$v4707\ := \$v4706\(0 to 3);
                \$v4705\ := \$v4706\(4 to 35);
                case \$v4707\ is
                when "0000" =>
                  \$12597\ := eclat_false;
                when "0001" =>
                  \$12613_j\ := \$v4705\(0 to 31);
                  \$12597\ := eclat_eq(\$12611_i\ & \$12613_j\);
                when others =>
                  
                end case;
                \$v4703\ := \$12597\;
                if \$v4703\(0) = '1' then
                  \$v4701\ := \$12587\(36 to 71);
                  \$v4702\ := \$v4701\(0 to 3);
                  \$v4694\ := \$v4701\(4 to 35);
                  case \$v4702\ is
                  when "0001" =>
                    \$12605_i\ := \$v4694\(0 to 31);
                    \$v4696\ := \$12588\(36 to 71);
                    \$v4697\ := \$v4696\(0 to 3);
                    \$v4695\ := \$v4696\(4 to 35);
                    case \$v4697\ is
                    when "0000" =>
                      \$12598\ := eclat_false;
                    when "0001" =>
                      \$12607_j\ := \$v4695\(0 to 31);
                      \$12598\ := eclat_eq(\$12605_i\ & \$12607_j\);
                    when others =>
                      
                    end case;
                    \$v4693\ := \$12598\;
                    if \$v4693\(0) = '1' then
                      \$v4691\ := \$12587\(72 to 107);
                      \$v4692\ := \$v4691\(0 to 3);
                      \$v4684\ := \$v4691\(4 to 35);
                      case \$v4692\ is
                      when "0001" =>
                        \$12599_i\ := \$v4684\(0 to 31);
                        \$v4686\ := \$12588\(72 to 107);
                        \$v4687\ := \$v4686\(0 to 3);
                        \$v4685\ := \$v4686\(4 to 35);
                        case \$v4687\ is
                        when "0000" =>
                          \$12552\ := eclat_false;
                        when "0001" =>
                          \$12601_j\ := \$v4685\(0 to 31);
                          \$12552\ := eclat_eq(\$12599_i\ & \$12601_j\);
                        when others =>
                          
                        end case;
                        \$v4678\ := \$$10702_brk_ptr_take\;
                        if \$v4678\(0) = '1' then
                          state_var7021 <= q_wait4677;
                        else
                          \$$10702_brk_ptr_take\(0) := '1';
                          \$$10702_brk_ptr\ <= 0;
                          state_var7021 <= pause_getI4675;
                        end if;
                      when "0000" =>
                        \$12602_i\ := \$v4684\(0 to 31);
                        \$v4689\ := \$12588\(72 to 107);
                        \$v4690\ := \$v4689\(0 to 3);
                        \$v4688\ := \$v4689\(4 to 35);
                        case \$v4690\ is
                        when "0001" =>
                          \$12552\ := eclat_false;
                        when "0000" =>
                          \$12604_j\ := \$v4688\(0 to 31);
                          \$12552\ := eclat_eq(\$12602_i\ & \$12604_j\);
                        when others =>
                          
                        end case;
                        \$v4678\ := \$$10702_brk_ptr_take\;
                        if \$v4678\(0) = '1' then
                          state_var7021 <= q_wait4677;
                        else
                          \$$10702_brk_ptr_take\(0) := '1';
                          \$$10702_brk_ptr\ <= 0;
                          state_var7021 <= pause_getI4675;
                        end if;
                      when others =>
                        
                      end case;
                    else
                      \$12552\ := eclat_false;
                      \$v4678\ := \$$10702_brk_ptr_take\;
                      if \$v4678\(0) = '1' then
                        state_var7021 <= q_wait4677;
                      else
                        \$$10702_brk_ptr_take\(0) := '1';
                        \$$10702_brk_ptr\ <= 0;
                        state_var7021 <= pause_getI4675;
                      end if;
                    end if;
                  when "0000" =>
                    \$12608_i\ := \$v4694\(0 to 31);
                    \$v4699\ := \$12588\(36 to 71);
                    \$v4700\ := \$v4699\(0 to 3);
                    \$v4698\ := \$v4699\(4 to 35);
                    case \$v4700\ is
                    when "0001" =>
                      \$12598\ := eclat_false;
                    when "0000" =>
                      \$12610_j\ := \$v4698\(0 to 31);
                      \$12598\ := eclat_eq(\$12608_i\ & \$12610_j\);
                    when others =>
                      
                    end case;
                    \$v4693\ := \$12598\;
                    if \$v4693\(0) = '1' then
                      \$v4691\ := \$12587\(72 to 107);
                      \$v4692\ := \$v4691\(0 to 3);
                      \$v4684\ := \$v4691\(4 to 35);
                      case \$v4692\ is
                      when "0001" =>
                        \$12599_i\ := \$v4684\(0 to 31);
                        \$v4686\ := \$12588\(72 to 107);
                        \$v4687\ := \$v4686\(0 to 3);
                        \$v4685\ := \$v4686\(4 to 35);
                        case \$v4687\ is
                        when "0000" =>
                          \$12552\ := eclat_false;
                        when "0001" =>
                          \$12601_j\ := \$v4685\(0 to 31);
                          \$12552\ := eclat_eq(\$12599_i\ & \$12601_j\);
                        when others =>
                          
                        end case;
                        \$v4678\ := \$$10702_brk_ptr_take\;
                        if \$v4678\(0) = '1' then
                          state_var7021 <= q_wait4677;
                        else
                          \$$10702_brk_ptr_take\(0) := '1';
                          \$$10702_brk_ptr\ <= 0;
                          state_var7021 <= pause_getI4675;
                        end if;
                      when "0000" =>
                        \$12602_i\ := \$v4684\(0 to 31);
                        \$v4689\ := \$12588\(72 to 107);
                        \$v4690\ := \$v4689\(0 to 3);
                        \$v4688\ := \$v4689\(4 to 35);
                        case \$v4690\ is
                        when "0001" =>
                          \$12552\ := eclat_false;
                        when "0000" =>
                          \$12604_j\ := \$v4688\(0 to 31);
                          \$12552\ := eclat_eq(\$12602_i\ & \$12604_j\);
                        when others =>
                          
                        end case;
                        \$v4678\ := \$$10702_brk_ptr_take\;
                        if \$v4678\(0) = '1' then
                          state_var7021 <= q_wait4677;
                        else
                          \$$10702_brk_ptr_take\(0) := '1';
                          \$$10702_brk_ptr\ <= 0;
                          state_var7021 <= pause_getI4675;
                        end if;
                      when others =>
                        
                      end case;
                    else
                      \$12552\ := eclat_false;
                      \$v4678\ := \$$10702_brk_ptr_take\;
                      if \$v4678\(0) = '1' then
                        state_var7021 <= q_wait4677;
                      else
                        \$$10702_brk_ptr_take\(0) := '1';
                        \$$10702_brk_ptr\ <= 0;
                        state_var7021 <= pause_getI4675;
                      end if;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$12552\ := eclat_false;
                  \$v4678\ := \$$10702_brk_ptr_take\;
                  if \$v4678\(0) = '1' then
                    state_var7021 <= q_wait4677;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI4675;
                  end if;
                end if;
              when "0000" =>
                \$12614_i\ := \$v4704\(0 to 31);
                \$v4709\ := \$12588\(0 to 35);
                \$v4710\ := \$v4709\(0 to 3);
                \$v4708\ := \$v4709\(4 to 35);
                case \$v4710\ is
                when "0001" =>
                  \$12597\ := eclat_false;
                when "0000" =>
                  \$12616_j\ := \$v4708\(0 to 31);
                  \$12597\ := eclat_eq(\$12614_i\ & \$12616_j\);
                when others =>
                  
                end case;
                \$v4703\ := \$12597\;
                if \$v4703\(0) = '1' then
                  \$v4701\ := \$12587\(36 to 71);
                  \$v4702\ := \$v4701\(0 to 3);
                  \$v4694\ := \$v4701\(4 to 35);
                  case \$v4702\ is
                  when "0001" =>
                    \$12605_i\ := \$v4694\(0 to 31);
                    \$v4696\ := \$12588\(36 to 71);
                    \$v4697\ := \$v4696\(0 to 3);
                    \$v4695\ := \$v4696\(4 to 35);
                    case \$v4697\ is
                    when "0000" =>
                      \$12598\ := eclat_false;
                    when "0001" =>
                      \$12607_j\ := \$v4695\(0 to 31);
                      \$12598\ := eclat_eq(\$12605_i\ & \$12607_j\);
                    when others =>
                      
                    end case;
                    \$v4693\ := \$12598\;
                    if \$v4693\(0) = '1' then
                      \$v4691\ := \$12587\(72 to 107);
                      \$v4692\ := \$v4691\(0 to 3);
                      \$v4684\ := \$v4691\(4 to 35);
                      case \$v4692\ is
                      when "0001" =>
                        \$12599_i\ := \$v4684\(0 to 31);
                        \$v4686\ := \$12588\(72 to 107);
                        \$v4687\ := \$v4686\(0 to 3);
                        \$v4685\ := \$v4686\(4 to 35);
                        case \$v4687\ is
                        when "0000" =>
                          \$12552\ := eclat_false;
                        when "0001" =>
                          \$12601_j\ := \$v4685\(0 to 31);
                          \$12552\ := eclat_eq(\$12599_i\ & \$12601_j\);
                        when others =>
                          
                        end case;
                        \$v4678\ := \$$10702_brk_ptr_take\;
                        if \$v4678\(0) = '1' then
                          state_var7021 <= q_wait4677;
                        else
                          \$$10702_brk_ptr_take\(0) := '1';
                          \$$10702_brk_ptr\ <= 0;
                          state_var7021 <= pause_getI4675;
                        end if;
                      when "0000" =>
                        \$12602_i\ := \$v4684\(0 to 31);
                        \$v4689\ := \$12588\(72 to 107);
                        \$v4690\ := \$v4689\(0 to 3);
                        \$v4688\ := \$v4689\(4 to 35);
                        case \$v4690\ is
                        when "0001" =>
                          \$12552\ := eclat_false;
                        when "0000" =>
                          \$12604_j\ := \$v4688\(0 to 31);
                          \$12552\ := eclat_eq(\$12602_i\ & \$12604_j\);
                        when others =>
                          
                        end case;
                        \$v4678\ := \$$10702_brk_ptr_take\;
                        if \$v4678\(0) = '1' then
                          state_var7021 <= q_wait4677;
                        else
                          \$$10702_brk_ptr_take\(0) := '1';
                          \$$10702_brk_ptr\ <= 0;
                          state_var7021 <= pause_getI4675;
                        end if;
                      when others =>
                        
                      end case;
                    else
                      \$12552\ := eclat_false;
                      \$v4678\ := \$$10702_brk_ptr_take\;
                      if \$v4678\(0) = '1' then
                        state_var7021 <= q_wait4677;
                      else
                        \$$10702_brk_ptr_take\(0) := '1';
                        \$$10702_brk_ptr\ <= 0;
                        state_var7021 <= pause_getI4675;
                      end if;
                    end if;
                  when "0000" =>
                    \$12608_i\ := \$v4694\(0 to 31);
                    \$v4699\ := \$12588\(36 to 71);
                    \$v4700\ := \$v4699\(0 to 3);
                    \$v4698\ := \$v4699\(4 to 35);
                    case \$v4700\ is
                    when "0001" =>
                      \$12598\ := eclat_false;
                    when "0000" =>
                      \$12610_j\ := \$v4698\(0 to 31);
                      \$12598\ := eclat_eq(\$12608_i\ & \$12610_j\);
                    when others =>
                      
                    end case;
                    \$v4693\ := \$12598\;
                    if \$v4693\(0) = '1' then
                      \$v4691\ := \$12587\(72 to 107);
                      \$v4692\ := \$v4691\(0 to 3);
                      \$v4684\ := \$v4691\(4 to 35);
                      case \$v4692\ is
                      when "0001" =>
                        \$12599_i\ := \$v4684\(0 to 31);
                        \$v4686\ := \$12588\(72 to 107);
                        \$v4687\ := \$v4686\(0 to 3);
                        \$v4685\ := \$v4686\(4 to 35);
                        case \$v4687\ is
                        when "0000" =>
                          \$12552\ := eclat_false;
                        when "0001" =>
                          \$12601_j\ := \$v4685\(0 to 31);
                          \$12552\ := eclat_eq(\$12599_i\ & \$12601_j\);
                        when others =>
                          
                        end case;
                        \$v4678\ := \$$10702_brk_ptr_take\;
                        if \$v4678\(0) = '1' then
                          state_var7021 <= q_wait4677;
                        else
                          \$$10702_brk_ptr_take\(0) := '1';
                          \$$10702_brk_ptr\ <= 0;
                          state_var7021 <= pause_getI4675;
                        end if;
                      when "0000" =>
                        \$12602_i\ := \$v4684\(0 to 31);
                        \$v4689\ := \$12588\(72 to 107);
                        \$v4690\ := \$v4689\(0 to 3);
                        \$v4688\ := \$v4689\(4 to 35);
                        case \$v4690\ is
                        when "0001" =>
                          \$12552\ := eclat_false;
                        when "0000" =>
                          \$12604_j\ := \$v4688\(0 to 31);
                          \$12552\ := eclat_eq(\$12602_i\ & \$12604_j\);
                        when others =>
                          
                        end case;
                        \$v4678\ := \$$10702_brk_ptr_take\;
                        if \$v4678\(0) = '1' then
                          state_var7021 <= q_wait4677;
                        else
                          \$$10702_brk_ptr_take\(0) := '1';
                          \$$10702_brk_ptr\ <= 0;
                          state_var7021 <= pause_getI4675;
                        end if;
                      when others =>
                        
                      end case;
                    else
                      \$12552\ := eclat_false;
                      \$v4678\ := \$$10702_brk_ptr_take\;
                      if \$v4678\(0) = '1' then
                        state_var7021 <= q_wait4677;
                      else
                        \$$10702_brk_ptr_take\(0) := '1';
                        \$$10702_brk_ptr\ <= 0;
                        state_var7021 <= pause_getI4675;
                      end if;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$12552\ := eclat_false;
                  \$v4678\ := \$$10702_brk_ptr_take\;
                  if \$v4678\(0) = '1' then
                    state_var7021 <= q_wait4677;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI4675;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII4722 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12587\ := \$$10696_ram_value\;
              \$v4718\ := \$12543_x\;
              \$v4719\ := \$v4718\(0 to 3);
              \$v4713\ := \$v4718\(4 to 35);
              case \$v4719\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12621_forever3163219\;
              when "0000" =>
                \$12629_i\ := \$v4713\(0 to 31);
                \$v4717\ := \$$10696_ram_ptr_take\;
                if \$v4717\(0) = '1' then
                  state_var7021 <= q_wait4716;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$12629_i\));
                  state_var7021 <= pause_getI4714;
                end if;
              when others =>
                
              end case;
            when pause_getII4739 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12546\ := \$$10696_ram_value\;
              \$v4736\ := \$12546\(36 to 71);
              \$v4737\ := \$v4736\(0 to 3);
              \$v4735\ := \$v4736\(4 to 35);
              case \$v4737\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12648_forever3163221\;
              when "0000" =>
                \$12656_i\ := \$v4735\(0 to 31);
                \$12550\ := \$12656_i\;
                \$v4734\ := \$$10697_stack_ptr_take\;
                if \$v4734\(0) = '1' then
                  state_var7021 <= q_wait4733;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12550\;
                  state_var7021 <= pause_setI4731;
                end if;
              when others =>
                
              end case;
            when pause_getII4743 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12545\ := \$$10697_stack_value\;
              \$v4741\ := \$$10696_ram_ptr_take\;
              if \$v4741\(0) = '1' then
                state_var7021 <= q_wait4740;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12545\));
                state_var7021 <= pause_getI4738;
              end if;
            when pause_getII4754 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12538\ := \$$10696_ram_value\;
              \$v4751\ := \$12538\(36 to 71);
              \$v4752\ := \$v4751\(0 to 3);
              \$v4750\ := \$v4751\(4 to 35);
              case \$v4752\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12662_forever3163222\;
              when "0000" =>
                \$12670_i\ := \$v4750\(0 to 31);
                \$12542\ := \$12670_i\;
                \$v4749\ := \$$10697_stack_ptr_take\;
                if \$v4749\(0) = '1' then
                  state_var7021 <= q_wait4748;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12542\;
                  state_var7021 <= pause_setI4746;
                end if;
              when others =>
                
              end case;
            when pause_getII4758 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12537\ := \$$10697_stack_value\;
              \$v4756\ := \$$10696_ram_ptr_take\;
              if \$v4756\(0) = '1' then
                state_var7021 <= q_wait4755;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12537\));
                state_var7021 <= pause_getI4753;
              end if;
            when pause_getII4767 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12694\ := \$$10697_stack_value\;
              \$v4765\ := \$$10696_ram_ptr_take\;
              if \$v4765\(0) = '1' then
                state_var7021 <= q_wait4764;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4761\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12694\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12687\ & "0000" & \$12692\ & "0001" & \$v4761\;
                state_var7021 <= pause_setI4762;
              end if;
            when pause_getII4775 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12692\ := \$$10697_stack_value\;
              \$v4773\ := \$$10697_stack_ptr_take\;
              if \$v4773\(0) = '1' then
                state_var7021 <= q_wait4772;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12691_i\;
                state_var7021 <= pause_setI4770;
              end if;
            when pause_getII4779 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12691_i\ := \$$10702_brk_value\;
              \$v4777\ := \$$10697_stack_ptr_take\;
              if \$v4777\(0) = '1' then
                state_var7021 <= q_wait4776;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4774;
              end if;
            when pause_getII4783 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12691_i\ := \$$10702_brk_value\;
              \$v4777\ := \$$10697_stack_ptr_take\;
              if \$v4777\(0) = '1' then
                state_var7021 <= q_wait4776;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4774;
              end if;
            when pause_getII4791 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12699\ := \$$10702_brk_value\;
              \$v4789\ := \$$10702_brk_ptr_take\;
              if \$v4789\(0) = '1' then
                state_var7021 <= q_wait4788;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12699\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4786;
              end if;
            when pause_getII4796 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12690\ := \$$10695_limit_value\;
              \$v4794\ := eclat_eq(\$12689\ & eclat_sub(\$12690\ & X"0000000" & X"1"));
              if \$v4794\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12707_forever3163223\;
              else
                \$v4793\ := \$$10702_brk_ptr_take\;
                if \$v4793\(0) = '1' then
                  state_var7021 <= q_wait4792;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4790;
                end if;
              end if;
            when pause_getII4800 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12689\ := \$$10702_brk_value\;
              \$v4798\ := \$$10695_limit_ptr_take\;
              if \$v4798\(0) = '1' then
                state_var7021 <= q_wait4797;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4795;
              end if;
            when pause_getII4819 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12681\ := \$$10696_ram_value\;
              \$v4816\ := \$12681\(36 to 71);
              \$v4817\ := \$v4816\(0 to 3);
              \$v4815\ := \$v4816\(4 to 35);
              case \$v4817\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12747_forever3163226\;
              when "0000" =>
                \$12755_i\ := \$v4815\(0 to 31);
                \$12685\ := \$12755_i\;
                \$v4814\ := \$$10697_stack_ptr_take\;
                if \$v4814\(0) = '1' then
                  state_var7021 <= q_wait4813;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12685\;
                  state_var7021 <= pause_setI4811;
                end if;
              when others =>
                
              end case;
            when pause_getII4823 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12680\ := \$$10697_stack_value\;
              \$v4821\ := \$$10696_ram_ptr_take\;
              if \$v4821\(0) = '1' then
                state_var7021 <= q_wait4820;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12680\));
                state_var7021 <= pause_getI4818;
              end if;
            when pause_getII4834 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12673\ := \$$10696_ram_value\;
              \$v4831\ := \$12673\(36 to 71);
              \$v4832\ := \$v4831\(0 to 3);
              \$v4830\ := \$v4831\(4 to 35);
              case \$v4832\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12761_forever3163227\;
              when "0000" =>
                \$12769_i\ := \$v4830\(0 to 31);
                \$12677\ := \$12769_i\;
                \$v4829\ := \$$10697_stack_ptr_take\;
                if \$v4829\(0) = '1' then
                  state_var7021 <= q_wait4828;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12677\;
                  state_var7021 <= pause_setI4826;
                end if;
              when others =>
                
              end case;
            when pause_getII4838 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12672\ := \$$10697_stack_value\;
              \$v4836\ := \$$10696_ram_ptr_take\;
              if \$v4836\(0) = '1' then
                state_var7021 <= q_wait4835;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12672\));
                state_var7021 <= pause_getI4833;
              end if;
            when pause_getII4847 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12793\ := \$$10697_stack_value\;
              \$v4845\ := \$$10696_ram_ptr_take\;
              if \$v4845\(0) = '1' then
                state_var7021 <= q_wait4844;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4841\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12793\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12786\ & "0000" & \$12791\ & "0001" & \$v4841\;
                state_var7021 <= pause_setI4842;
              end if;
            when pause_getII4855 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12791\ := \$$10697_stack_value\;
              \$v4853\ := \$$10697_stack_ptr_take\;
              if \$v4853\(0) = '1' then
                state_var7021 <= q_wait4852;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12790_i\;
                state_var7021 <= pause_setI4850;
              end if;
            when pause_getII4859 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12790_i\ := \$$10702_brk_value\;
              \$v4857\ := \$$10697_stack_ptr_take\;
              if \$v4857\(0) = '1' then
                state_var7021 <= q_wait4856;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4854;
              end if;
            when pause_getII4863 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12790_i\ := \$$10702_brk_value\;
              \$v4857\ := \$$10697_stack_ptr_take\;
              if \$v4857\(0) = '1' then
                state_var7021 <= q_wait4856;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4854;
              end if;
            when pause_getII4871 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12798\ := \$$10702_brk_value\;
              \$v4869\ := \$$10702_brk_ptr_take\;
              if \$v4869\(0) = '1' then
                state_var7021 <= q_wait4868;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12798\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4866;
              end if;
            when pause_getII4876 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12789\ := \$$10695_limit_value\;
              \$v4874\ := eclat_eq(\$12788\ & eclat_sub(\$12789\ & X"0000000" & X"1"));
              if \$v4874\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12806_forever3163228\;
              else
                \$v4873\ := \$$10702_brk_ptr_take\;
                if \$v4873\(0) = '1' then
                  state_var7021 <= q_wait4872;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4870;
                end if;
              end if;
            when pause_getII4880 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12788\ := \$$10702_brk_value\;
              \$v4878\ := \$$10695_limit_ptr_take\;
              if \$v4878\(0) = '1' then
                state_var7021 <= q_wait4877;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4875;
              end if;
            when pause_getII4898 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12780\ := \$$10696_ram_value\;
              \$v4895\ := \$12780\(36 to 71);
              \$v4896\ := \$v4895\(0 to 3);
              \$v4894\ := \$v4895\(4 to 35);
              case \$v4896\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12847_forever3163231\;
              when "0000" =>
                \$12855_i\ := \$v4894\(0 to 31);
                \$12784\ := \$12855_i\;
                \$v4893\ := \$$10697_stack_ptr_take\;
                if \$v4893\(0) = '1' then
                  state_var7021 <= q_wait4892;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12784\;
                  state_var7021 <= pause_setI4890;
                end if;
              when others =>
                
              end case;
            when pause_getII4902 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12779\ := \$$10697_stack_value\;
              \$v4900\ := \$$10696_ram_ptr_take\;
              if \$v4900\(0) = '1' then
                state_var7021 <= q_wait4899;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12779\));
                state_var7021 <= pause_getI4897;
              end if;
            when pause_getII4913 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12772\ := \$$10696_ram_value\;
              \$v4910\ := \$12772\(36 to 71);
              \$v4911\ := \$v4910\(0 to 3);
              \$v4909\ := \$v4910\(4 to 35);
              case \$v4911\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12861_forever3163232\;
              when "0000" =>
                \$12869_i\ := \$v4909\(0 to 31);
                \$12776\ := \$12869_i\;
                \$v4908\ := \$$10697_stack_ptr_take\;
                if \$v4908\(0) = '1' then
                  state_var7021 <= q_wait4907;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12776\;
                  state_var7021 <= pause_setI4905;
                end if;
              when others =>
                
              end case;
            when pause_getII4917 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12771\ := \$$10697_stack_value\;
              \$v4915\ := \$$10696_ram_ptr_take\;
              if \$v4915\(0) = '1' then
                state_var7021 <= q_wait4914;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12771\));
                state_var7021 <= pause_getI4912;
              end if;
            when pause_getII4926 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12893\ := \$$10697_stack_value\;
              \$v4924\ := \$$10696_ram_ptr_take\;
              if \$v4924\(0) = '1' then
                state_var7021 <= q_wait4923;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4920\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12893\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12886\ & "0000" & \$12891\ & "0001" & \$v4920\;
                state_var7021 <= pause_setI4921;
              end if;
            when pause_getII4934 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12891\ := \$$10697_stack_value\;
              \$v4932\ := \$$10697_stack_ptr_take\;
              if \$v4932\(0) = '1' then
                state_var7021 <= q_wait4931;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12890_i\;
                state_var7021 <= pause_setI4929;
              end if;
            when pause_getII4938 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12890_i\ := \$$10702_brk_value\;
              \$v4936\ := \$$10697_stack_ptr_take\;
              if \$v4936\(0) = '1' then
                state_var7021 <= q_wait4935;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4933;
              end if;
            when pause_getII4942 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12890_i\ := \$$10702_brk_value\;
              \$v4936\ := \$$10697_stack_ptr_take\;
              if \$v4936\(0) = '1' then
                state_var7021 <= q_wait4935;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4933;
              end if;
            when pause_getII4950 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12898\ := \$$10702_brk_value\;
              \$v4948\ := \$$10702_brk_ptr_take\;
              if \$v4948\(0) = '1' then
                state_var7021 <= q_wait4947;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12898\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4945;
              end if;
            when pause_getII4955 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12889\ := \$$10695_limit_value\;
              \$v4953\ := eclat_eq(\$12888\ & eclat_sub(\$12889\ & X"0000000" & X"1"));
              if \$v4953\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12906_forever3163233\;
              else
                \$v4952\ := \$$10702_brk_ptr_take\;
                if \$v4952\(0) = '1' then
                  state_var7021 <= q_wait4951;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4949;
                end if;
              end if;
            when pause_getII4959 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12888\ := \$$10702_brk_value\;
              \$v4957\ := \$$10695_limit_ptr_take\;
              if \$v4957\(0) = '1' then
                state_var7021 <= q_wait4956;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4954;
              end if;
            when pause_getII4977 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12880\ := \$$10696_ram_value\;
              \$v4974\ := \$12880\(36 to 71);
              \$v4975\ := \$v4974\(0 to 3);
              \$v4973\ := \$v4974\(4 to 35);
              case \$v4975\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12947_forever3163236\;
              when "0000" =>
                \$12955_i\ := \$v4973\(0 to 31);
                \$12884\ := \$12955_i\;
                \$v4972\ := \$$10697_stack_ptr_take\;
                if \$v4972\(0) = '1' then
                  state_var7021 <= q_wait4971;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12884\;
                  state_var7021 <= pause_setI4969;
                end if;
              when others =>
                
              end case;
            when pause_getII4981 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12879\ := \$$10697_stack_value\;
              \$v4979\ := \$$10696_ram_ptr_take\;
              if \$v4979\(0) = '1' then
                state_var7021 <= q_wait4978;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12879\));
                state_var7021 <= pause_getI4976;
              end if;
            when pause_getII4992 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12872\ := \$$10696_ram_value\;
              \$v4989\ := \$12872\(36 to 71);
              \$v4990\ := \$v4989\(0 to 3);
              \$v4988\ := \$v4989\(4 to 35);
              case \$v4990\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12961_forever3163237\;
              when "0000" =>
                \$12969_i\ := \$v4988\(0 to 31);
                \$12876\ := \$12969_i\;
                \$v4987\ := \$$10697_stack_ptr_take\;
                if \$v4987\(0) = '1' then
                  state_var7021 <= q_wait4986;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12876\;
                  state_var7021 <= pause_setI4984;
                end if;
              when others =>
                
              end case;
            when pause_getII4996 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12871\ := \$$10697_stack_value\;
              \$v4994\ := \$$10696_ram_ptr_take\;
              if \$v4994\(0) = '1' then
                state_var7021 <= q_wait4993;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12871\));
                state_var7021 <= pause_getI4991;
              end if;
            when pause_getII5005 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12993\ := \$$10697_stack_value\;
              \$v5003\ := \$$10696_ram_ptr_take\;
              if \$v5003\(0) = '1' then
                state_var7021 <= q_wait5002;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4999\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12993\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12986\ & "0000" & \$12991\ & "0001" & \$v4999\;
                state_var7021 <= pause_setI5000;
              end if;
            when pause_getII5013 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12991\ := \$$10697_stack_value\;
              \$v5011\ := \$$10697_stack_ptr_take\;
              if \$v5011\(0) = '1' then
                state_var7021 <= q_wait5010;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12990_i\;
                state_var7021 <= pause_setI5008;
              end if;
            when pause_getII5017 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12990_i\ := \$$10702_brk_value\;
              \$v5015\ := \$$10697_stack_ptr_take\;
              if \$v5015\(0) = '1' then
                state_var7021 <= q_wait5014;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5012;
              end if;
            when pause_getII5021 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12990_i\ := \$$10702_brk_value\;
              \$v5015\ := \$$10697_stack_ptr_take\;
              if \$v5015\(0) = '1' then
                state_var7021 <= q_wait5014;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5012;
              end if;
            when pause_getII5029 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12998\ := \$$10702_brk_value\;
              \$v5027\ := \$$10702_brk_ptr_take\;
              if \$v5027\(0) = '1' then
                state_var7021 <= q_wait5026;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12998\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5024;
              end if;
            when pause_getII5034 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$12989\ := \$$10695_limit_value\;
              \$v5032\ := eclat_eq(\$12988\ & eclat_sub(\$12989\ & X"0000000" & X"1"));
              if \$v5032\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13006_forever3163238\;
              else
                \$v5031\ := \$$10702_brk_ptr_take\;
                if \$v5031\(0) = '1' then
                  state_var7021 <= q_wait5030;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5028;
                end if;
              end if;
            when pause_getII5038 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$12988\ := \$$10702_brk_value\;
              \$v5036\ := \$$10695_limit_ptr_take\;
              if \$v5036\(0) = '1' then
                state_var7021 <= q_wait5035;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5033;
              end if;
            when pause_getII5056 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12980\ := \$$10696_ram_value\;
              \$v5053\ := \$12980\(36 to 71);
              \$v5054\ := \$v5053\(0 to 3);
              \$v5052\ := \$v5053\(4 to 35);
              case \$v5054\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13047_forever3163241\;
              when "0000" =>
                \$13055_i\ := \$v5052\(0 to 31);
                \$12984\ := \$13055_i\;
                \$v5051\ := \$$10697_stack_ptr_take\;
                if \$v5051\(0) = '1' then
                  state_var7021 <= q_wait5050;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12984\;
                  state_var7021 <= pause_setI5048;
                end if;
              when others =>
                
              end case;
            when pause_getII5060 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12979\ := \$$10697_stack_value\;
              \$v5058\ := \$$10696_ram_ptr_take\;
              if \$v5058\(0) = '1' then
                state_var7021 <= q_wait5057;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12979\));
                state_var7021 <= pause_getI5055;
              end if;
            when pause_getII5071 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$12972\ := \$$10696_ram_value\;
              \$v5068\ := \$12972\(36 to 71);
              \$v5069\ := \$v5068\(0 to 3);
              \$v5067\ := \$v5068\(4 to 35);
              case \$v5069\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13061_forever3163242\;
              when "0000" =>
                \$13069_i\ := \$v5067\(0 to 31);
                \$12976\ := \$13069_i\;
                \$v5066\ := \$$10697_stack_ptr_take\;
                if \$v5066\(0) = '1' then
                  state_var7021 <= q_wait5065;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$12976\;
                  state_var7021 <= pause_setI5063;
                end if;
              when others =>
                
              end case;
            when pause_getII5075 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12971\ := \$$10697_stack_value\;
              \$v5073\ := \$$10696_ram_ptr_take\;
              if \$v5073\(0) = '1' then
                state_var7021 <= q_wait5072;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12971\));
                state_var7021 <= pause_getI5070;
              end if;
            when pause_getII5084 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13093\ := \$$10697_stack_value\;
              \$v5082\ := \$$10696_ram_ptr_take\;
              if \$v5082\(0) = '1' then
                state_var7021 <= q_wait5081;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5078\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13093\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13086\ & "0000" & \$13091\ & "0001" & \$v5078\;
                state_var7021 <= pause_setI5079;
              end if;
            when pause_getII5092 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13091\ := \$$10697_stack_value\;
              \$v5090\ := \$$10697_stack_ptr_take\;
              if \$v5090\(0) = '1' then
                state_var7021 <= q_wait5089;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13090_i\;
                state_var7021 <= pause_setI5087;
              end if;
            when pause_getII5096 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13090_i\ := \$$10702_brk_value\;
              \$v5094\ := \$$10697_stack_ptr_take\;
              if \$v5094\(0) = '1' then
                state_var7021 <= q_wait5093;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5091;
              end if;
            when pause_getII5100 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13090_i\ := \$$10702_brk_value\;
              \$v5094\ := \$$10697_stack_ptr_take\;
              if \$v5094\(0) = '1' then
                state_var7021 <= q_wait5093;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5091;
              end if;
            when pause_getII5108 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13098\ := \$$10702_brk_value\;
              \$v5106\ := \$$10702_brk_ptr_take\;
              if \$v5106\(0) = '1' then
                state_var7021 <= q_wait5105;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13098\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5103;
              end if;
            when pause_getII5113 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$13089\ := \$$10695_limit_value\;
              \$v5111\ := eclat_eq(\$13088\ & eclat_sub(\$13089\ & X"0000000" & X"1"));
              if \$v5111\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13106_forever3163243\;
              else
                \$v5110\ := \$$10702_brk_ptr_take\;
                if \$v5110\(0) = '1' then
                  state_var7021 <= q_wait5109;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5107;
                end if;
              end if;
            when pause_getII5117 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13088\ := \$$10702_brk_value\;
              \$v5115\ := \$$10695_limit_ptr_take\;
              if \$v5115\(0) = '1' then
                state_var7021 <= q_wait5114;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5112;
              end if;
            when pause_getII5135 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13080\ := \$$10696_ram_value\;
              \$v5132\ := \$13080\(36 to 71);
              \$v5133\ := \$v5132\(0 to 3);
              \$v5131\ := \$v5132\(4 to 35);
              case \$v5133\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13147_forever3163246\;
              when "0000" =>
                \$13155_i\ := \$v5131\(0 to 31);
                \$13084\ := \$13155_i\;
                \$v5130\ := \$$10697_stack_ptr_take\;
                if \$v5130\(0) = '1' then
                  state_var7021 <= q_wait5129;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$13084\;
                  state_var7021 <= pause_setI5127;
                end if;
              when others =>
                
              end case;
            when pause_getII5139 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13079\ := \$$10697_stack_value\;
              \$v5137\ := \$$10696_ram_ptr_take\;
              if \$v5137\(0) = '1' then
                state_var7021 <= q_wait5136;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13079\));
                state_var7021 <= pause_getI5134;
              end if;
            when pause_getII5150 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13072\ := \$$10696_ram_value\;
              \$v5147\ := \$13072\(36 to 71);
              \$v5148\ := \$v5147\(0 to 3);
              \$v5146\ := \$v5147\(4 to 35);
              case \$v5148\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13161_forever3163247\;
              when "0000" =>
                \$13169_i\ := \$v5146\(0 to 31);
                \$13076\ := \$13169_i\;
                \$v5145\ := \$$10697_stack_ptr_take\;
                if \$v5145\(0) = '1' then
                  state_var7021 <= q_wait5144;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$13076\;
                  state_var7021 <= pause_setI5142;
                end if;
              when others =>
                
              end case;
            when pause_getII5154 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13071\ := \$$10697_stack_value\;
              \$v5152\ := \$$10696_ram_ptr_take\;
              if \$v5152\(0) = '1' then
                state_var7021 <= q_wait5151;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13071\));
                state_var7021 <= pause_getI5149;
              end if;
            when pause_getII5163 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13181\ := \$$10697_stack_value\;
              \$v5161\ := \$$10696_ram_ptr_take\;
              if \$v5161\(0) = '1' then
                state_var7021 <= q_wait5160;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5157\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13181\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13174\ & "0000" & \$13179\ & "0001" & \$v5157\;
                state_var7021 <= pause_setI5158;
              end if;
            when pause_getII5171 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13179\ := \$$10697_stack_value\;
              \$v5169\ := \$$10697_stack_ptr_take\;
              if \$v5169\(0) = '1' then
                state_var7021 <= q_wait5168;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13178_i\;
                state_var7021 <= pause_setI5166;
              end if;
            when pause_getII5175 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13178_i\ := \$$10702_brk_value\;
              \$v5173\ := \$$10697_stack_ptr_take\;
              if \$v5173\(0) = '1' then
                state_var7021 <= q_wait5172;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5170;
              end if;
            when pause_getII5179 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13178_i\ := \$$10702_brk_value\;
              \$v5173\ := \$$10697_stack_ptr_take\;
              if \$v5173\(0) = '1' then
                state_var7021 <= q_wait5172;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5170;
              end if;
            when pause_getII5187 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13186\ := \$$10702_brk_value\;
              \$v5185\ := \$$10702_brk_ptr_take\;
              if \$v5185\(0) = '1' then
                state_var7021 <= q_wait5184;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13186\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5182;
              end if;
            when pause_getII5192 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$13177\ := \$$10695_limit_value\;
              \$v5190\ := eclat_eq(\$13176\ & eclat_sub(\$13177\ & X"0000000" & X"1"));
              if \$v5190\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13194_forever3163248\;
              else
                \$v5189\ := \$$10702_brk_ptr_take\;
                if \$v5189\(0) = '1' then
                  state_var7021 <= q_wait5188;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5186;
                end if;
              end if;
            when pause_getII5196 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13176\ := \$$10702_brk_value\;
              \$v5194\ := \$$10695_limit_ptr_take\;
              if \$v5194\(0) = '1' then
                state_var7021 <= q_wait5193;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5191;
              end if;
            when pause_getII5205 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13229\ := \$$10697_stack_value\;
              \$v5203\ := \$$10696_ram_ptr_take\;
              if \$v5203\(0) = '1' then
                state_var7021 <= q_wait5202;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5199\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13229\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13222\ & "0000" & \$13227\ & "0001" & \$v5199\;
                state_var7021 <= pause_setI5200;
              end if;
            when pause_getII5213 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13227\ := \$$10697_stack_value\;
              \$v5211\ := \$$10697_stack_ptr_take\;
              if \$v5211\(0) = '1' then
                state_var7021 <= q_wait5210;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13226_i\;
                state_var7021 <= pause_setI5208;
              end if;
            when pause_getII5217 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13226_i\ := \$$10702_brk_value\;
              \$v5215\ := \$$10697_stack_ptr_take\;
              if \$v5215\(0) = '1' then
                state_var7021 <= q_wait5214;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5212;
              end if;
            when pause_getII5221 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13226_i\ := \$$10702_brk_value\;
              \$v5215\ := \$$10697_stack_ptr_take\;
              if \$v5215\(0) = '1' then
                state_var7021 <= q_wait5214;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5212;
              end if;
            when pause_getII5229 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13234\ := \$$10702_brk_value\;
              \$v5227\ := \$$10702_brk_ptr_take\;
              if \$v5227\(0) = '1' then
                state_var7021 <= q_wait5226;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13234\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5224;
              end if;
            when pause_getII5234 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$13225\ := \$$10695_limit_value\;
              \$v5232\ := eclat_eq(\$13224\ & eclat_sub(\$13225\ & X"0000000" & X"1"));
              if \$v5232\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13242_forever3163250\;
              else
                \$v5231\ := \$$10702_brk_ptr_take\;
                if \$v5231\(0) = '1' then
                  state_var7021 <= q_wait5230;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5228;
                end if;
              end if;
            when pause_getII5238 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13224\ := \$$10702_brk_value\;
              \$v5236\ := \$$10695_limit_ptr_take\;
              if \$v5236\(0) = '1' then
                state_var7021 <= q_wait5235;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5233;
              end if;
            when pause_getII5252 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13216\ := \$$10696_ram_value\;
              \$v5249\ := \$13216\(36 to 71);
              \$v5250\ := \$v5249\(0 to 3);
              \$v5248\ := \$v5249\(4 to 35);
              case \$v5250\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13270_forever3163252\;
              when "0000" =>
                \$13278_i\ := \$v5248\(0 to 31);
                \$13220\ := \$13278_i\;
                \$v5247\ := \$$10697_stack_ptr_take\;
                if \$v5247\(0) = '1' then
                  state_var7021 <= q_wait5246;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$13220\;
                  state_var7021 <= pause_setI5244;
                end if;
              when others =>
                
              end case;
            when pause_getII5256 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13215\ := \$$10697_stack_value\;
              \$v5254\ := \$$10696_ram_ptr_take\;
              if \$v5254\(0) = '1' then
                state_var7021 <= q_wait5253;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13215\));
                state_var7021 <= pause_getI5251;
              end if;
            when pause_getII5264 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10819\ := \$$10696_ram_value\;
              \$v5260\ := \$10819\(0 to 35);
              \$v5261\ := \$v5260\(0 to 3);
              \$v3369\ := \$v5260\(4 to 35);
              case \$v5261\ is
              when "0000" =>
                \$v3629\ := \$$10702_brk_ptr_take\;
                if \$v3629\(0) = '1' then
                  state_var7021 <= q_wait3628;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI3626;
                end if;
              when "0001" =>
                \$11321_i\ := \$v3369\(0 to 31);
                \$v5259\ := \$11321_i\;
                case \$v5259\ is
                when X"0000000" & X"0" =>
                  \$v3847\ := \$$10697_stack_ptr_take\;
                  if \$v3847\(0) = '1' then
                    state_var7021 <= q_wait3846;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI3844;
                  end if;
                when X"0000000" & X"1" =>
                  \$v3904\ := \$$10697_stack_ptr_take\;
                  if \$v3904\(0) = '1' then
                    state_var7021 <= q_wait3903;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI3901;
                  end if;
                when X"0000000" & X"2" =>
                  \$v3919\ := \$$10697_stack_ptr_take\;
                  if \$v3919\(0) = '1' then
                    state_var7021 <= q_wait3918;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI3916;
                  end if;
                when X"0000000" & X"3" =>
                  \$v3991\ := \$$10697_stack_ptr_take\;
                  if \$v3991\(0) = '1' then
                    state_var7021 <= q_wait3990;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI3988;
                  end if;
                when X"0000000" & X"4" =>
                  \$v4101\ := \$$10697_stack_ptr_take\;
                  if \$v4101\(0) = '1' then
                    state_var7021 <= q_wait4100;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4098;
                  end if;
                when X"0000000" & X"5" =>
                  \$v4163\ := \$$10697_stack_ptr_take\;
                  if \$v4163\(0) = '1' then
                    state_var7021 <= q_wait4162;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4160;
                  end if;
                when X"0000000" & X"6" =>
                  \$v4227\ := \$$10697_stack_ptr_take\;
                  if \$v4227\(0) = '1' then
                    state_var7021 <= q_wait4226;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4224;
                  end if;
                when X"0000000" & X"7" =>
                  \$v4291\ := \$$10697_stack_ptr_take\;
                  if \$v4291\(0) = '1' then
                    state_var7021 <= q_wait4290;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4288;
                  end if;
                when X"0000000" & X"8" =>
                  \$v4355\ := \$$10697_stack_ptr_take\;
                  if \$v4355\(0) = '1' then
                    state_var7021 <= q_wait4354;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4352;
                  end if;
                when X"0000000" & X"9" =>
                  \$v4448\ := \$$10697_stack_ptr_take\;
                  if \$v4448\(0) = '1' then
                    state_var7021 <= q_wait4447;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4445;
                  end if;
                when X"0000000" & X"a" =>
                  \$v4541\ := \$$10697_stack_ptr_take\;
                  if \$v4541\(0) = '1' then
                    state_var7021 <= q_wait4540;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4538;
                  end if;
                when X"0000000" & X"b" =>
                  \$v4634\ := \$$10697_stack_ptr_take\;
                  if \$v4634\(0) = '1' then
                    state_var7021 <= q_wait4633;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4631;
                  end if;
                when X"0000000" & X"c" =>
                  \$v4760\ := \$$10697_stack_ptr_take\;
                  if \$v4760\(0) = '1' then
                    state_var7021 <= q_wait4759;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4757;
                  end if;
                when X"0000000" & X"d" =>
                  \$v4840\ := \$$10697_stack_ptr_take\;
                  if \$v4840\(0) = '1' then
                    state_var7021 <= q_wait4839;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4837;
                  end if;
                when X"0000000" & X"e" =>
                  \$v4919\ := \$$10697_stack_ptr_take\;
                  if \$v4919\(0) = '1' then
                    state_var7021 <= q_wait4918;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4916;
                  end if;
                when X"0000000" & X"f" =>
                  \$v4998\ := \$$10697_stack_ptr_take\;
                  if \$v4998\(0) = '1' then
                    state_var7021 <= q_wait4997;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI4995;
                  end if;
                when X"000000" & X"10" =>
                  \$v5077\ := \$$10697_stack_ptr_take\;
                  if \$v5077\(0) = '1' then
                    state_var7021 <= q_wait5076;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI5074;
                  end if;
                when X"000000" & X"11" =>
                  \$v5156\ := \$$10697_stack_ptr_take\;
                  if \$v5156\(0) = '1' then
                    state_var7021 <= q_wait5155;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI5153;
                  end if;
                when X"000000" & X"12" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("get_char is not available"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13206_forever3163249\;
                when X"000000" & X"13" =>
                  \$v5258\ := \$$10697_stack_ptr_take\;
                  if \$v5258\(0) = '1' then
                    state_var7021 <= q_wait5257;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI5255;
                  end if;
                when others =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("invalid primitive identifier"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$11525_forever3163173\;
                end case;
              when others =>
                
              end case;
            when pause_getII5272 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13296\ := \$$10696_ram_value\;
              \$10818_proc\ := \$13296\(0 to 35);
              \$v5267\ := \$10818_proc\;
              \$v5268\ := \$v5267\(0 to 3);
              \$v5262\ := \$v5267\(4 to 35);
              case \$v5268\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13283_forever3163253\;
              when "0000" =>
                \$13291_i\ := \$v5262\(0 to 31);
                \$v5266\ := \$$10696_ram_ptr_take\;
                if \$v5266\(0) = '1' then
                  state_var7021 <= q_wait5265;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13291_i\));
                  state_var7021 <= pause_getI5263;
                end if;
              when others =>
                
              end case;
            when pause_getII5279 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13327\ := \$$10696_ram_value\;
              \$13318_list_tail2653256_arg\ := \$13327\(36 to 71) & eclat_sub(\$13318_list_tail2653256_arg\(36 to 67) & X"0000000" & X"1") & eclat_unit;
              state_var7021 <= \$13318_list_tail2653256\;
            when pause_getII5286 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13294\ := \$$10697_stack_value\;
              \$13318_list_tail2653256_arg\ := "0000" & \$13294\ & \$13292_i\ & eclat_unit;
              state_var7021 <= \$13318_list_tail2653256\;
            when pause_getII5291 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13351\ := \$$10696_ram_value\;
              \$10818_proc\ := \$13351\(0 to 35);
              \$v5267\ := \$10818_proc\;
              \$v5268\ := \$v5267\(0 to 3);
              \$v5262\ := \$v5267\(4 to 35);
              case \$v5268\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13283_forever3163253\;
              when "0000" =>
                \$13291_i\ := \$v5262\(0 to 31);
                \$v5266\ := \$$10696_ram_ptr_take\;
                if \$v5266\(0) = '1' then
                  state_var7021 <= q_wait5265;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13291_i\));
                  state_var7021 <= pause_getI5263;
                end if;
              when others =>
                
              end case;
            when pause_getII5300 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10814\ := \$$10696_ram_value\;
              \$v5296\ := \$10814\(36 to 71);
              \$v5297\ := \$v5296\(0 to 3);
              \$v5269\ := \$v5296\(4 to 35);
              case \$v5297\ is
              when "0001" =>
                \$13292_i\ := \$v5269\(0 to 31);
                \$v5288\ := \$$10697_stack_ptr_take\;
                if \$v5288\(0) = '1' then
                  state_var7021 <= q_wait5287;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI5285;
                end if;
              when "0000" =>
                \$v5294\ := \$10814\(36 to 71);
                \$v5295\ := \$v5294\(0 to 3);
                \$v5289\ := \$v5294\(4 to 35);
                case \$v5295\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13360_forever3163257\;
                when "0000" =>
                  \$13368_i\ := \$v5289\(0 to 31);
                  \$v5293\ := \$$10696_ram_ptr_take\;
                  if \$v5293\(0) = '1' then
                    state_var7021 <= q_wait5292;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$13368_i\));
                    state_var7021 <= pause_getI5290;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII5306 =>
              \$$10700_pc_ptr_take\(0) := '0';
              \$10813\ := \$$10700_pc_value\;
              \$v5303\ := "0000" & \$10813\;
              \$v5304\ := \$v5303\(0 to 3);
              \$v5298\ := \$v5303\(4 to 35);
              case \$v5304\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13374_forever3163258\;
              when "0000" =>
                \$13382_i\ := \$v5298\(0 to 31);
                \$v5302\ := \$$10696_ram_ptr_take\;
                if \$v5302\(0) = '1' then
                  state_var7021 <= q_wait5301;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13382_i\));
                  state_var7021 <= pause_getI5299;
                end if;
              when others =>
                
              end case;
            when pause_getII5311 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10811\ := \$$10702_brk_value\;
              \$v5309\ := eclat_lt(eclat_sub(\$10810\ & \$10811\) & X"000000" & X"32");
              if \$v5309\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13388_forever3163259\;
              else
                \$v5308\ := \$$10700_pc_ptr_take\;
                if \$v5308\(0) = '1' then
                  state_var7021 <= q_wait5307;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI5305;
                end if;
              end if;
            when pause_getII5315 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$10810\ := \$$10695_limit_value\;
              \$v5313\ := \$$10702_brk_ptr_take\;
              if \$v5313\(0) = '1' then
                state_var7021 <= q_wait5312;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5310;
              end if;
            when pause_getII5327 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13409\ := \$$10696_ram_value\;
              \$v5323\ := \$13409\(72 to 107);
              \$v5324\ := \$v5323\(0 to 3);
              \$v5322\ := \$v5323\(4 to 35);
              case \$v5324\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13420_forever3163260\;
              when "0000" =>
                \$13428_i\ := \$v5322\(0 to 31);
                \$13415\ := \$13428_i\;
                \$v5321\ := \$$10700_pc_ptr_take\;
                if \$v5321\(0) = '1' then
                  state_var7021 <= q_wait5320;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr_write\ <= 0;
                  \$$10700_pc_write_request\ <= '1';
                  \$$10700_pc_write\ <= \$13415\;
                  state_var7021 <= pause_setI5318;
                end if;
              when others =>
                
              end case;
            when pause_getII5333 =>
              \$$10700_pc_ptr_take\(0) := '0';
              \$13408\ := \$$10700_pc_value\;
              \$v5330\ := "0000" & \$13408\;
              \$v5331\ := \$v5330\(0 to 3);
              \$v5325\ := \$v5330\(4 to 35);
              case \$v5331\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13434_forever3163261\;
              when "0000" =>
                \$13442_i\ := \$v5325\(0 to 31);
                \$v5329\ := \$$10696_ram_ptr_take\;
                if \$v5329\(0) = '1' then
                  state_var7021 <= q_wait5328;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13442_i\));
                  state_var7021 <= pause_getI5326;
                end if;
              when others =>
                
              end case;
            when pause_getII5344 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13461\ := \$$10696_ram_value\;
              \$v5341\ := \$$10696_ram_ptr_take\;
              if \$v5341\(0) = '1' then
                state_var7021 <= q_wait5340;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13459_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13405\ & \$13460\(36 to 71) & \$13461\(72 to 107);
                state_var7021 <= pause_setI5338;
              end if;
            when pause_getII5351 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13460\ := \$$10696_ram_value\;
              \$v5347\ := \$13446\;
              \$v5348\ := \$v5347\(0 to 3);
              \$v5342\ := \$v5347\(4 to 35);
              case \$v5348\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13474_forever3163263\;
              when "0000" =>
                \$13482_i\ := \$v5342\(0 to 31);
                \$v5346\ := \$$10696_ram_ptr_take\;
                if \$v5346\(0) = '1' then
                  state_var7021 <= q_wait5345;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13482_i\));
                  state_var7021 <= pause_getI5343;
                end if;
              when others =>
                
              end case;
            when pause_getII5360 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13509\ := \$$10696_ram_value\;
              \$13500_list_tail2653266_arg\ := \$13509\(36 to 71) & eclat_sub(\$13500_list_tail2653266_arg\(36 to 67) & X"0000000" & X"1") & eclat_unit;
              state_var7021 <= \$13500_list_tail2653266\;
            when pause_getII5367 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13445\ := \$$10697_stack_value\;
              \$13500_list_tail2653266_arg\ := "0000" & \$13445\ & \$13443_i\ & eclat_unit;
              state_var7021 <= \$13500_list_tail2653266\;
            when pause_getII5377 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13547\ := \$$10696_ram_value\;
              \$v5374\ := \$$10696_ram_ptr_take\;
              if \$v5374\(0) = '1' then
                state_var7021 <= q_wait5373;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13545_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13405\ & \$13546\(36 to 71) & \$13547\(72 to 107);
                state_var7021 <= pause_setI5371;
              end if;
            when pause_getII5384 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13546\ := \$$10696_ram_value\;
              \$v5380\ := \$10793\(36 to 71);
              \$v5381\ := \$v5380\(0 to 3);
              \$v5375\ := \$v5380\(4 to 35);
              case \$v5381\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13560_forever3163268\;
              when "0000" =>
                \$13568_i\ := \$v5375\(0 to 31);
                \$v5379\ := \$$10696_ram_ptr_take\;
                if \$v5379\(0) = '1' then
                  state_var7021 <= q_wait5378;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13568_i\));
                  state_var7021 <= pause_getI5376;
                end if;
              when others =>
                
              end case;
            when pause_getII5401 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13400\ := \$$10696_ram_value\;
              \$v5398\ := \$13400\(36 to 71);
              \$v5399\ := \$v5398\(0 to 3);
              \$v5397\ := \$v5398\(4 to 35);
              case \$v5399\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13587_forever3163270\;
              when "0000" =>
                \$13595_i\ := \$v5397\(0 to 31);
                \$13404\ := \$13595_i\;
                \$v5396\ := \$$10697_stack_ptr_take\;
                if \$v5396\(0) = '1' then
                  state_var7021 <= q_wait5395;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$13404\;
                  state_var7021 <= pause_setI5393;
                end if;
              when others =>
                
              end case;
            when pause_getII5405 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13399\ := \$$10697_stack_value\;
              \$v5403\ := \$$10696_ram_ptr_take\;
              if \$v5403\(0) = '1' then
                state_var7021 <= q_wait5402;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13399\));
                state_var7021 <= pause_getI5400;
              end if;
            when pause_getII5417 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13607\ := \$$10696_ram_value\;
              \$v5413\ := \$13607\(72 to 107);
              \$v5414\ := \$v5413\(0 to 3);
              \$v5412\ := \$v5413\(4 to 35);
              case \$v5414\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13618_forever3163271\;
              when "0000" =>
                \$13626_i\ := \$v5412\(0 to 31);
                \$13613\ := \$13626_i\;
                \$v5411\ := \$$10700_pc_ptr_take\;
                if \$v5411\(0) = '1' then
                  state_var7021 <= q_wait5410;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr_write\ <= 0;
                  \$$10700_pc_write_request\ <= '1';
                  \$$10700_pc_write\ <= \$13613\;
                  state_var7021 <= pause_setI5408;
                end if;
              when others =>
                
              end case;
            when pause_getII5423 =>
              \$$10700_pc_ptr_take\(0) := '0';
              \$13606\ := \$$10700_pc_value\;
              \$v5420\ := "0000" & \$13606\;
              \$v5421\ := \$v5420\(0 to 3);
              \$v5415\ := \$v5420\(4 to 35);
              case \$v5421\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13632_forever3163272\;
              when "0000" =>
                \$13640_i\ := \$v5415\(0 to 31);
                \$v5419\ := \$$10696_ram_ptr_take\;
                if \$v5419\(0) = '1' then
                  state_var7021 <= q_wait5418;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13640_i\));
                  state_var7021 <= pause_getI5416;
                end if;
              when others =>
                
              end case;
            when pause_getII5432 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13603\ := \$$10697_stack_value\;
              \$v5430\ := \$$10696_ram_ptr_take\;
              if \$v5430\(0) = '1' then
                state_var7021 <= q_wait5429;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5426\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13603\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13596_v\ & "0000" & \$13601\ & "0001" & \$v5426\;
                state_var7021 <= pause_setI5427;
              end if;
            when pause_getII5440 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13601\ := \$$10697_stack_value\;
              \$v5438\ := \$$10697_stack_ptr_take\;
              if \$v5438\(0) = '1' then
                state_var7021 <= q_wait5437;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13600_i\;
                state_var7021 <= pause_setI5435;
              end if;
            when pause_getII5444 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13600_i\ := \$$10702_brk_value\;
              \$v5442\ := \$$10697_stack_ptr_take\;
              if \$v5442\(0) = '1' then
                state_var7021 <= q_wait5441;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5439;
              end if;
            when pause_getII5448 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13600_i\ := \$$10702_brk_value\;
              \$v5442\ := \$$10697_stack_ptr_take\;
              if \$v5442\(0) = '1' then
                state_var7021 <= q_wait5441;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5439;
              end if;
            when pause_getII5456 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13645\ := \$$10702_brk_value\;
              \$v5454\ := \$$10702_brk_ptr_take\;
              if \$v5454\(0) = '1' then
                state_var7021 <= q_wait5453;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13645\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5451;
              end if;
            when pause_getII5461 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$13599\ := \$$10695_limit_value\;
              \$v5459\ := eclat_eq(\$13598\ & eclat_sub(\$13599\ & X"0000000" & X"1"));
              if \$v5459\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13653_forever3163273\;
              else
                \$v5458\ := \$$10702_brk_ptr_take\;
                if \$v5458\(0) = '1' then
                  state_var7021 <= q_wait5457;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5455;
                end if;
              end if;
            when pause_getII5465 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13598\ := \$$10702_brk_value\;
              \$v5463\ := \$$10695_limit_ptr_take\;
              if \$v5463\(0) = '1' then
                state_var7021 <= q_wait5462;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5460;
              end if;
            when pause_getII5471 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13667\ := \$$10696_ram_value\;
              \$13596_v\ := \$13667\(0 to 35);
              \$v5467\ := \$$10702_brk_ptr_take\;
              if \$v5467\(0) = '1' then
                state_var7021 <= q_wait5466;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5464;
              end if;
            when pause_getII5478 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13698\ := \$$10696_ram_value\;
              \$13689_list_tail2653276_arg\ := \$13698\(36 to 71) & eclat_sub(\$13689_list_tail2653276_arg\(36 to 67) & X"0000000" & X"1") & eclat_unit;
              state_var7021 <= \$13689_list_tail2653276\;
            when pause_getII5485 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13665\ := \$$10697_stack_value\;
              \$13689_list_tail2653276_arg\ := "0000" & \$13665\ & \$13663_i\ & eclat_unit;
              state_var7021 <= \$13689_list_tail2653276\;
            when pause_getII5490 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13722\ := \$$10696_ram_value\;
              \$13596_v\ := \$13722\(0 to 35);
              \$v5467\ := \$$10702_brk_ptr_take\;
              if \$v5467\(0) = '1' then
                state_var7021 <= q_wait5466;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5464;
              end if;
            when pause_getII5506 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13750\ := \$$10696_ram_value\;
              \$v5502\ := \$13750\(72 to 107);
              \$v5503\ := \$v5502\(0 to 3);
              \$v5501\ := \$v5502\(4 to 35);
              case \$v5503\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13761_forever3163278\;
              when "0000" =>
                \$13769_i\ := \$v5501\(0 to 31);
                \$13756\ := \$13769_i\;
                \$v5500\ := \$$10700_pc_ptr_take\;
                if \$v5500\(0) = '1' then
                  state_var7021 <= q_wait5499;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr_write\ <= 0;
                  \$$10700_pc_write_request\ <= '1';
                  \$$10700_pc_write\ <= \$13756\;
                  state_var7021 <= pause_setI5497;
                end if;
              when others =>
                
              end case;
            when pause_getII5512 =>
              \$$10700_pc_ptr_take\(0) := '0';
              \$13749\ := \$$10700_pc_value\;
              \$v5509\ := "0000" & \$13749\;
              \$v5510\ := \$v5509\(0 to 3);
              \$v5504\ := \$v5509\(4 to 35);
              case \$v5510\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13775_forever3163279\;
              when "0000" =>
                \$13783_i\ := \$v5504\(0 to 31);
                \$v5508\ := \$$10696_ram_ptr_take\;
                if \$v5508\(0) = '1' then
                  state_var7021 <= q_wait5507;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13783_i\));
                  state_var7021 <= pause_getI5505;
                end if;
              when others =>
                
              end case;
            when pause_getII5521 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13746\ := \$$10697_stack_value\;
              \$v5519\ := \$$10696_ram_ptr_take\;
              if \$v5519\(0) = '1' then
                state_var7021 <= q_wait5518;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5515\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13746\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$10793\(36 to 71) & "0000" & \$13744\ & "0001" & \$v5515\;
                state_var7021 <= pause_setI5516;
              end if;
            when pause_getII5529 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13744\ := \$$10697_stack_value\;
              \$v5527\ := \$$10697_stack_ptr_take\;
              if \$v5527\(0) = '1' then
                state_var7021 <= q_wait5526;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13743_i\;
                state_var7021 <= pause_setI5524;
              end if;
            when pause_getII5533 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13743_i\ := \$$10702_brk_value\;
              \$v5531\ := \$$10697_stack_ptr_take\;
              if \$v5531\(0) = '1' then
                state_var7021 <= q_wait5530;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5528;
              end if;
            when pause_getII5537 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13743_i\ := \$$10702_brk_value\;
              \$v5531\ := \$$10697_stack_ptr_take\;
              if \$v5531\(0) = '1' then
                state_var7021 <= q_wait5530;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5528;
              end if;
            when pause_getII5545 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13788\ := \$$10702_brk_value\;
              \$v5543\ := \$$10702_brk_ptr_take\;
              if \$v5543\(0) = '1' then
                state_var7021 <= q_wait5542;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13788\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5540;
              end if;
            when pause_getII5550 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$13742\ := \$$10695_limit_value\;
              \$v5548\ := eclat_eq(\$13741\ & eclat_sub(\$13742\ & X"0000000" & X"1"));
              if \$v5548\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13796_forever3163280\;
              else
                \$v5547\ := \$$10702_brk_ptr_take\;
                if \$v5547\(0) = '1' then
                  state_var7021 <= q_wait5546;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5544;
                end if;
              end if;
            when pause_getII5554 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13741\ := \$$10702_brk_value\;
              \$v5552\ := \$$10695_limit_ptr_take\;
              if \$v5552\(0) = '1' then
                state_var7021 <= q_wait5551;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5549;
              end if;
            when pause_getII5566 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13832\ := \$$10696_ram_value\;
              \$v5562\ := \$13832\(72 to 107);
              \$v5563\ := \$v5562\(0 to 3);
              \$v5561\ := \$v5562\(4 to 35);
              case \$v5563\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13842_forever3163282\;
              when "0000" =>
                \$13850_i\ := \$v5561\(0 to 31);
                \$13837\ := \$13850_i\;
                \$v5560\ := \$$10700_pc_ptr_take\;
                if \$v5560\(0) = '1' then
                  state_var7021 <= q_wait5559;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr_write\ <= 0;
                  \$$10700_pc_write_request\ <= '1';
                  \$$10700_pc_write\ <= \$13837\;
                  state_var7021 <= pause_setI5557;
                end if;
              when others =>
                
              end case;
            when pause_getII5572 =>
              \$$10700_pc_ptr_take\(0) := '0';
              \$13831\ := \$$10700_pc_value\;
              \$v5569\ := "0000" & \$13831\;
              \$v5570\ := \$v5569\(0 to 3);
              \$v5564\ := \$v5569\(4 to 35);
              case \$v5570\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13856_forever3163283\;
              when "0000" =>
                \$13864_i\ := \$v5564\(0 to 31);
                \$v5568\ := \$$10696_ram_ptr_take\;
                if \$v5568\(0) = '1' then
                  state_var7021 <= q_wait5567;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13864_i\));
                  state_var7021 <= pause_getI5565;
                end if;
              when others =>
                
              end case;
            when pause_getII5602 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13808\ := \$$10696_ram_value\;
              \$v5599\ := \$13808\(36 to 71);
              \$v5600\ := \$v5599\(0 to 3);
              \$v5598\ := \$v5599\(4 to 35);
              case \$v5600\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13878_forever3163284\;
              when "0000" =>
                \$13886_i\ := \$v5598\(0 to 31);
                \$13812\ := \$13886_i\;
                \$v5597\ := \$$10697_stack_ptr_take\;
                if \$v5597\(0) = '1' then
                  state_var7021 <= q_wait5596;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$13812\;
                  state_var7021 <= pause_setI5594;
                end if;
              when others =>
                
              end case;
            when pause_getII5606 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13807\ := \$$10697_stack_value\;
              \$v5604\ := \$$10696_ram_ptr_take\;
              if \$v5604\(0) = '1' then
                state_var7021 <= q_wait5603;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13807\));
                state_var7021 <= pause_getI5601;
              end if;
            when pause_getII5614 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10793\ := \$$10696_ram_value\;
              \$v5610\ := \$10793\(0 to 35);
              \$v5611\ := \$v5610\(0 to 3);
              \$v3368\ := \$v5610\(4 to 35);
              case \$v5611\ is
              when "0001" =>
                \$10797_i\ := \$v3368\(0 to 31);
                \$v5609\ := \$10797_i\;
                case \$v5609\ is
                when X"0000000" & X"0" =>
                  \$v5317\ := \$$10695_limit_ptr_take\;
                  if \$v5317\(0) = '1' then
                    state_var7021 <= q_wait5316;
                  else
                    \$$10695_limit_ptr_take\(0) := '1';
                    \$$10695_limit_ptr\ <= 0;
                    state_var7021 <= pause_getI5314;
                  end if;
                when X"0000000" & X"1" =>
                  \$v5407\ := \$$10697_stack_ptr_take\;
                  if \$v5407\(0) = '1' then
                    state_var7021 <= q_wait5406;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI5404;
                  end if;
                when X"0000000" & X"2" =>
                  \$v5495\ := \$10793\(36 to 71);
                  \$v5496\ := \$v5495\(0 to 3);
                  \$v5468\ := \$v5495\(4 to 35);
                  case \$v5496\ is
                  when "0001" =>
                    \$13663_i\ := \$v5468\(0 to 31);
                    \$v5487\ := \$$10697_stack_ptr_take\;
                    if \$v5487\(0) = '1' then
                      state_var7021 <= q_wait5486;
                    else
                      \$$10697_stack_ptr_take\(0) := '1';
                      \$$10697_stack_ptr\ <= 0;
                      state_var7021 <= pause_getI5484;
                    end if;
                  when "0000" =>
                    \$v5493\ := \$10793\(36 to 71);
                    \$v5494\ := \$v5493\(0 to 3);
                    \$v5488\ := \$v5493\(4 to 35);
                    case \$v5494\ is
                    when "0001" =>
                      eclat_print_string(of_string("Fatal error : "));
                      
                      eclat_print_string(of_string("can't get_rib"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var7021 <= \$13731_forever3163277\;
                    when "0000" =>
                      \$13739_i\ := \$v5488\(0 to 31);
                      \$v5492\ := \$$10696_ram_ptr_take\;
                      if \$v5492\(0) = '1' then
                        state_var7021 <= q_wait5491;
                      else
                        \$$10696_ram_ptr_take\(0) := '1';
                        \$$10696_ram_ptr\ <= to_integer(unsigned(\$13739_i\));
                        state_var7021 <= pause_getI5489;
                      end if;
                    when others =>
                      
                    end case;
                  when others =>
                    
                  end case;
                when X"0000000" & X"3" =>
                  \$v5556\ := \$$10702_brk_ptr_take\;
                  if \$v5556\(0) = '1' then
                    state_var7021 <= q_wait5555;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI5553;
                  end if;
                when X"0000000" & X"4" =>
                  \$v5608\ := \$$10697_stack_ptr_take\;
                  if \$v5608\(0) = '1' then
                    state_var7021 <= q_wait5607;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI5605;
                  end if;
                when X"0000000" & X"5" =>
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("HALT!"));
                  
                  \$10778_run286_result\ := eclat_unit;
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$10704_forever290\;
                when others =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("not implemented yet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$10801_forever3163135\;
                end case;
              when others =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented yet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13892_forever3163134\;
              end case;
            when pause_getII5620 =>
              \$$10700_pc_ptr_take\(0) := '0';
              \$10792\ := \$$10700_pc_value\;
              \$v5617\ := "0000" & \$10792\;
              \$v5618\ := \$v5617\(0 to 3);
              \$v5612\ := \$v5617\(4 to 35);
              case \$v5618\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13905_forever3163285\;
              when "0000" =>
                \$13913_i\ := \$v5612\(0 to 31);
                \$v5616\ := \$$10696_ram_ptr_take\;
                if \$v5616\(0) = '1' then
                  state_var7021 <= q_wait5615;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13913_i\));
                  state_var7021 <= pause_getI5613;
                end if;
              when others =>
                
              end case;
            when pause_getII5641 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10767_j\ := \$$10702_brk_value\;
              \$v5639\ := \$$10696_ram_ptr_take\;
              if \$v5639\(0) = '1' then
                state_var7021 <= q_wait5638;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5633\ := X"0000000" & X"5";
                \$v5634\ := X"0000000" & X"0";
                \$v5635\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10763_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5633\ & "0001" & \$v5634\ & "0001" & \$v5635\;
                state_var7021 <= pause_setI5636;
              end if;
            when pause_getII5645 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10767_j\ := \$$10702_brk_value\;
              \$v5639\ := \$$10696_ram_ptr_take\;
              if \$v5639\(0) = '1' then
                state_var7021 <= q_wait5638;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5633\ := X"0000000" & X"5";
                \$v5634\ := X"0000000" & X"0";
                \$v5635\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10763_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5633\ & "0001" & \$v5634\ & "0001" & \$v5635\;
                state_var7021 <= pause_setI5636;
              end if;
            when pause_getII5653 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13923\ := \$$10702_brk_value\;
              \$v5651\ := \$$10702_brk_ptr_take\;
              if \$v5651\(0) = '1' then
                state_var7021 <= q_wait5650;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13923\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5648;
              end if;
            when pause_getII5658 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$10766\ := \$$10695_limit_value\;
              \$v5656\ := eclat_eq(\$10765\ & eclat_sub(\$10766\ & X"0000000" & X"1"));
              if \$v5656\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13931_forever3163286\;
              else
                \$v5655\ := \$$10702_brk_ptr_take\;
                if \$v5655\(0) = '1' then
                  state_var7021 <= q_wait5654;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5652;
                end if;
              end if;
            when pause_getII5662 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10765\ := \$$10702_brk_value\;
              \$v5660\ := \$$10695_limit_ptr_take\;
              if \$v5660\(0) = '1' then
                state_var7021 <= q_wait5659;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5657;
              end if;
            when pause_getII5666 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10763_i\ := \$$10702_brk_value\;
              \$v5664\ := \$$10702_brk_ptr_take\;
              if \$v5664\(0) = '1' then
                state_var7021 <= q_wait5663;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5661;
              end if;
            when pause_getII5670 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10763_i\ := \$$10702_brk_value\;
              \$v5664\ := \$$10702_brk_ptr_take\;
              if \$v5664\(0) = '1' then
                state_var7021 <= q_wait5663;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5661;
              end if;
            when pause_getII5678 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$13942\ := \$$10702_brk_value\;
              \$v5676\ := \$$10702_brk_ptr_take\;
              if \$v5676\(0) = '1' then
                state_var7021 <= q_wait5675;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13942\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5673;
              end if;
            when pause_getII5683 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$10762\ := \$$10695_limit_value\;
              \$v5681\ := eclat_eq(\$10761\ & eclat_sub(\$10762\ & X"0000000" & X"1"));
              if \$v5681\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13950_forever3163287\;
              else
                \$v5680\ := \$$10702_brk_ptr_take\;
                if \$v5680\(0) = '1' then
                  state_var7021 <= q_wait5679;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5677;
                end if;
              end if;
            when pause_getII5687 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10761\ := \$$10702_brk_value\;
              \$v5685\ := \$$10695_limit_ptr_take\;
              if \$v5685\(0) = '1' then
                state_var7021 <= q_wait5684;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5682;
              end if;
            when pause_getII5699 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$13967\ := \$$10696_ram_value\;
              \$v5695\ := \$13967\(36 to 71);
              \$v5696\ := \$v5695\(0 to 3);
              \$v5694\ := \$v5695\(4 to 35);
              case \$v5696\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13977_forever3163288\;
              when "0000" =>
                \$13985_i\ := \$v5694\(0 to 31);
                \$13972\ := \$13985_i\;
                \$v5693\ := \$$10699_symtbl_ptr_take\;
                if \$v5693\(0) = '1' then
                  state_var7021 <= q_wait5692;
                else
                  \$$10699_symtbl_ptr_take\(0) := '1';
                  \$$10699_symtbl_ptr_write\ <= 0;
                  \$$10699_symtbl_write_request\ <= '1';
                  \$$10699_symtbl_write\ <= \$13972\;
                  state_var7021 <= pause_setI5690;
                end if;
              when others =>
                
              end case;
            when pause_getII5705 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$13966\ := \$$10699_symtbl_value\;
              \$v5702\ := "0000" & \$13966\;
              \$v5703\ := \$v5702\(0 to 3);
              \$v5697\ := \$v5702\(4 to 35);
              case \$v5703\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13991_forever3163289\;
              when "0000" =>
                \$13999_i\ := \$v5697\(0 to 31);
                \$v5701\ := \$$10696_ram_ptr_take\;
                if \$v5701\(0) = '1' then
                  state_var7021 <= q_wait5700;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$13999_i\));
                  state_var7021 <= pause_getI5698;
                end if;
              when others =>
                
              end case;
            when pause_getII5716 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14022\ := \$$10696_ram_value\;
              \$v5713\ := \$$10696_ram_ptr_take\;
              if \$v5713\(0) = '1' then
                state_var7021 <= q_wait5712;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5709\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14012_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v5709\ & \$14017\(36 to 71) & \$14022\(72 to 107);
                state_var7021 <= pause_setI5710;
              end if;
            when pause_getII5723 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14017\ := \$$10696_ram_value\;
              \$v5719\ := \$10758\(0 to 35);
              \$v5720\ := \$v5719\(0 to 3);
              \$v5714\ := \$v5719\(4 to 35);
              case \$v5720\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14037_forever3163291\;
              when "0000" =>
                \$14045_i\ := \$v5714\(0 to 31);
                \$v5718\ := \$$10696_ram_ptr_take\;
                if \$v5718\(0) = '1' then
                  state_var7021 <= q_wait5717;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14045_i\));
                  state_var7021 <= pause_getI5715;
                end if;
              when others =>
                
              end case;
            when pause_getII5732 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10758\ := \$$10696_ram_value\;
              \$v5728\ := \$10758\(0 to 35);
              \$v5729\ := \$v5728\(0 to 3);
              \$v5708\ := \$v5728\(4 to 35);
              case \$v5729\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14004_forever3163290\;
              when "0000" =>
                \$14012_i\ := \$v5708\(0 to 31);
                \$v5726\ := \$10758\(0 to 35);
                \$v5727\ := \$v5726\(0 to 3);
                \$v5721\ := \$v5726\(4 to 35);
                case \$v5727\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14050_forever3163292\;
                when "0000" =>
                  \$14058_i\ := \$v5721\(0 to 31);
                  \$v5725\ := \$$10696_ram_ptr_take\;
                  if \$v5725\(0) = '1' then
                    state_var7021 <= q_wait5724;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14058_i\));
                    state_var7021 <= pause_getI5722;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII5738 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$10757\ := \$$10699_symtbl_value\;
              \$v5735\ := "0000" & \$10757\;
              \$v5736\ := \$v5735\(0 to 3);
              \$v5730\ := \$v5735\(4 to 35);
              case \$v5736\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14064_forever3163293\;
              when "0000" =>
                \$14072_i\ := \$v5730\(0 to 31);
                \$v5734\ := \$$10696_ram_ptr_take\;
                if \$v5734\(0) = '1' then
                  state_var7021 <= q_wait5733;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14072_i\));
                  state_var7021 <= pause_getI5731;
                end if;
              when others =>
                
              end case;
            when pause_getII5750 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14080\ := \$$10696_ram_value\;
              \$v5746\ := \$14080\(36 to 71);
              \$v5747\ := \$v5746\(0 to 3);
              \$v5745\ := \$v5746\(4 to 35);
              case \$v5747\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14090_forever3163294\;
              when "0000" =>
                \$14098_i\ := \$v5745\(0 to 31);
                \$14085\ := \$14098_i\;
                \$v5744\ := \$$10699_symtbl_ptr_take\;
                if \$v5744\(0) = '1' then
                  state_var7021 <= q_wait5743;
                else
                  \$$10699_symtbl_ptr_take\(0) := '1';
                  \$$10699_symtbl_ptr_write\ <= 0;
                  \$$10699_symtbl_write_request\ <= '1';
                  \$$10699_symtbl_write\ <= \$14085\;
                  state_var7021 <= pause_setI5741;
                end if;
              when others =>
                
              end case;
            when pause_getII5756 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$14079\ := \$$10699_symtbl_value\;
              \$v5753\ := "0000" & \$14079\;
              \$v5754\ := \$v5753\(0 to 3);
              \$v5748\ := \$v5753\(4 to 35);
              case \$v5754\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14104_forever3163295\;
              when "0000" =>
                \$14112_i\ := \$v5748\(0 to 31);
                \$v5752\ := \$$10696_ram_ptr_take\;
                if \$v5752\(0) = '1' then
                  state_var7021 <= q_wait5751;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14112_i\));
                  state_var7021 <= pause_getI5749;
                end if;
              when others =>
                
              end case;
            when pause_getII5767 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14135\ := \$$10696_ram_value\;
              \$v5764\ := \$$10696_ram_ptr_take\;
              if \$v5764\(0) = '1' then
                state_var7021 <= q_wait5763;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5760\ := X"0000000" & X"1";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14125_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v5760\ & \$14130\(36 to 71) & \$14135\(72 to 107);
                state_var7021 <= pause_setI5761;
              end if;
            when pause_getII5774 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14130\ := \$$10696_ram_value\;
              \$v5770\ := \$10754\(0 to 35);
              \$v5771\ := \$v5770\(0 to 3);
              \$v5765\ := \$v5770\(4 to 35);
              case \$v5771\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14150_forever3163297\;
              when "0000" =>
                \$14158_i\ := \$v5765\(0 to 31);
                \$v5769\ := \$$10696_ram_ptr_take\;
                if \$v5769\(0) = '1' then
                  state_var7021 <= q_wait5768;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14158_i\));
                  state_var7021 <= pause_getI5766;
                end if;
              when others =>
                
              end case;
            when pause_getII5783 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10754\ := \$$10696_ram_value\;
              \$v5779\ := \$10754\(0 to 35);
              \$v5780\ := \$v5779\(0 to 3);
              \$v5759\ := \$v5779\(4 to 35);
              case \$v5780\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14117_forever3163296\;
              when "0000" =>
                \$14125_i\ := \$v5759\(0 to 31);
                \$v5777\ := \$10754\(0 to 35);
                \$v5778\ := \$v5777\(0 to 3);
                \$v5772\ := \$v5777\(4 to 35);
                case \$v5778\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14163_forever3163298\;
                when "0000" =>
                  \$14171_i\ := \$v5772\(0 to 31);
                  \$v5776\ := \$$10696_ram_ptr_take\;
                  if \$v5776\(0) = '1' then
                    state_var7021 <= q_wait5775;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14171_i\));
                    state_var7021 <= pause_getI5773;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII5789 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$10753\ := \$$10699_symtbl_value\;
              \$v5786\ := "0000" & \$10753\;
              \$v5787\ := \$v5786\(0 to 3);
              \$v5781\ := \$v5786\(4 to 35);
              case \$v5787\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14177_forever3163299\;
              when "0000" =>
                \$14185_i\ := \$v5781\(0 to 31);
                \$v5785\ := \$$10696_ram_ptr_take\;
                if \$v5785\(0) = '1' then
                  state_var7021 <= q_wait5784;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14185_i\));
                  state_var7021 <= pause_getI5782;
                end if;
              when others =>
                
              end case;
            when pause_getII5801 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14193\ := \$$10696_ram_value\;
              \$v5797\ := \$14193\(36 to 71);
              \$v5798\ := \$v5797\(0 to 3);
              \$v5796\ := \$v5797\(4 to 35);
              case \$v5798\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14203_forever3163300\;
              when "0000" =>
                \$14211_i\ := \$v5796\(0 to 31);
                \$14198\ := \$14211_i\;
                \$v5795\ := \$$10699_symtbl_ptr_take\;
                if \$v5795\(0) = '1' then
                  state_var7021 <= q_wait5794;
                else
                  \$$10699_symtbl_ptr_take\(0) := '1';
                  \$$10699_symtbl_ptr_write\ <= 0;
                  \$$10699_symtbl_write_request\ <= '1';
                  \$$10699_symtbl_write\ <= \$14198\;
                  state_var7021 <= pause_setI5792;
                end if;
              when others =>
                
              end case;
            when pause_getII5807 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$14192\ := \$$10699_symtbl_value\;
              \$v5804\ := "0000" & \$14192\;
              \$v5805\ := \$v5804\(0 to 3);
              \$v5799\ := \$v5804\(4 to 35);
              case \$v5805\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14217_forever3163301\;
              when "0000" =>
                \$14225_i\ := \$v5799\(0 to 31);
                \$v5803\ := \$$10696_ram_ptr_take\;
                if \$v5803\(0) = '1' then
                  state_var7021 <= q_wait5802;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14225_i\));
                  state_var7021 <= pause_getI5800;
                end if;
              when others =>
                
              end case;
            when pause_getII5818 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14248\ := \$$10696_ram_value\;
              \$v5815\ := \$$10696_ram_ptr_take\;
              if \$v5815\(0) = '1' then
                state_var7021 <= q_wait5814;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5811\ := X"0000000" & X"2";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14238_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v5811\ & \$14243\(36 to 71) & \$14248\(72 to 107);
                state_var7021 <= pause_setI5812;
              end if;
            when pause_getII5825 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14243\ := \$$10696_ram_value\;
              \$v5821\ := \$10750\(0 to 35);
              \$v5822\ := \$v5821\(0 to 3);
              \$v5816\ := \$v5821\(4 to 35);
              case \$v5822\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14263_forever3163303\;
              when "0000" =>
                \$14271_i\ := \$v5816\(0 to 31);
                \$v5820\ := \$$10696_ram_ptr_take\;
                if \$v5820\(0) = '1' then
                  state_var7021 <= q_wait5819;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14271_i\));
                  state_var7021 <= pause_getI5817;
                end if;
              when others =>
                
              end case;
            when pause_getII5834 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10750\ := \$$10696_ram_value\;
              \$v5830\ := \$10750\(0 to 35);
              \$v5831\ := \$v5830\(0 to 3);
              \$v5810\ := \$v5830\(4 to 35);
              case \$v5831\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14230_forever3163302\;
              when "0000" =>
                \$14238_i\ := \$v5810\(0 to 31);
                \$v5828\ := \$10750\(0 to 35);
                \$v5829\ := \$v5828\(0 to 3);
                \$v5823\ := \$v5828\(4 to 35);
                case \$v5829\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14276_forever3163304\;
                when "0000" =>
                  \$14284_i\ := \$v5823\(0 to 31);
                  \$v5827\ := \$$10696_ram_ptr_take\;
                  if \$v5827\(0) = '1' then
                    state_var7021 <= q_wait5826;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14284_i\));
                    state_var7021 <= pause_getI5824;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII5840 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$10749\ := \$$10699_symtbl_value\;
              \$v5837\ := "0000" & \$10749\;
              \$v5838\ := \$v5837\(0 to 3);
              \$v5832\ := \$v5837\(4 to 35);
              case \$v5838\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14290_forever3163305\;
              when "0000" =>
                \$14298_i\ := \$v5832\(0 to 31);
                \$v5836\ := \$$10696_ram_ptr_take\;
                if \$v5836\(0) = '1' then
                  state_var7021 <= q_wait5835;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14298_i\));
                  state_var7021 <= pause_getI5833;
                end if;
              when others =>
                
              end case;
            when pause_getII5852 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14301\ := \$$10696_ram_value\;
              \$v5848\ := \$14301\(36 to 71);
              \$v5849\ := \$v5848\(0 to 3);
              \$v5847\ := \$v5848\(4 to 35);
              case \$v5849\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14311_forever3163306\;
              when "0000" =>
                \$14319_i\ := \$v5847\(0 to 31);
                \$14306\ := \$14319_i\;
                \$v5846\ := \$$10699_symtbl_ptr_take\;
                if \$v5846\(0) = '1' then
                  state_var7021 <= q_wait5845;
                else
                  \$$10699_symtbl_ptr_take\(0) := '1';
                  \$$10699_symtbl_ptr_write\ <= 0;
                  \$$10699_symtbl_write_request\ <= '1';
                  \$$10699_symtbl_write\ <= \$14306\;
                  state_var7021 <= pause_setI5843;
                end if;
              when others =>
                
              end case;
            when pause_getII5858 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$14300\ := \$$10699_symtbl_value\;
              \$v5855\ := "0000" & \$14300\;
              \$v5856\ := \$v5855\(0 to 3);
              \$v5850\ := \$v5855\(4 to 35);
              case \$v5856\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14325_forever3163307\;
              when "0000" =>
                \$14333_i\ := \$v5850\(0 to 31);
                \$v5854\ := \$$10696_ram_ptr_take\;
                if \$v5854\(0) = '1' then
                  state_var7021 <= q_wait5853;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14333_i\));
                  state_var7021 <= pause_getI5851;
                end if;
              when others =>
                
              end case;
            when pause_getII5868 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14356\ := \$$10696_ram_value\;
              \$v5865\ := \$$10696_ram_ptr_take\;
              if \$v5865\(0) = '1' then
                state_var7021 <= q_wait5864;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14346_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$10738_main_rib\ & \$14351\(36 to 71) & \$14356\(72 to 107);
                state_var7021 <= pause_setI5862;
              end if;
            when pause_getII5875 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14351\ := \$$10696_ram_value\;
              \$v5871\ := \$10741\(0 to 35);
              \$v5872\ := \$v5871\(0 to 3);
              \$v5866\ := \$v5871\(4 to 35);
              case \$v5872\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14369_forever3163309\;
              when "0000" =>
                \$14377_i\ := \$v5866\(0 to 31);
                \$v5870\ := \$$10696_ram_ptr_take\;
                if \$v5870\(0) = '1' then
                  state_var7021 <= q_wait5869;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14377_i\));
                  state_var7021 <= pause_getI5867;
                end if;
              when others =>
                
              end case;
            when pause_getII5884 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10741\ := \$$10696_ram_value\;
              \$v5880\ := \$10741\(0 to 35);
              \$v5881\ := \$v5880\(0 to 3);
              \$v5861\ := \$v5880\(4 to 35);
              case \$v5881\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14338_forever3163308\;
              when "0000" =>
                \$14346_i\ := \$v5861\(0 to 31);
                \$v5878\ := \$10741\(0 to 35);
                \$v5879\ := \$v5878\(0 to 3);
                \$v5873\ := \$v5878\(4 to 35);
                case \$v5879\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14382_forever3163310\;
                when "0000" =>
                  \$14390_i\ := \$v5873\(0 to 31);
                  \$v5877\ := \$$10696_ram_ptr_take\;
                  if \$v5877\(0) = '1' then
                    state_var7021 <= q_wait5876;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14390_i\));
                    state_var7021 <= pause_getI5874;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII5890 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$10740\ := \$$10699_symtbl_value\;
              \$v5887\ := "0000" & \$10740\;
              \$v5888\ := \$v5887\(0 to 3);
              \$v5882\ := \$v5887\(4 to 35);
              case \$v5888\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14396_forever3163311\;
              when "0000" =>
                \$14404_i\ := \$v5882\(0 to 31);
                \$v5886\ := \$$10696_ram_ptr_take\;
                if \$v5886\(0) = '1' then
                  state_var7021 <= q_wait5885;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14404_i\));
                  state_var7021 <= pause_getI5883;
                end if;
              when others =>
                
              end case;
            when pause_getII5894 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14409\ := \$$10698_heap_value\;
              \$10738_main_rib\ := "0000" & \$14409\;
              \$v5892\ := \$$10699_symtbl_ptr_take\;
              if \$v5892\(0) = '1' then
                state_var7021 <= q_wait5891;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5889;
              end if;
            when pause_getII5904 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14407\ := \$$10698_heap_value\;
              \$v5902\ := \$$10696_ram_ptr_take\;
              if \$v5902\(0) = '1' then
                state_var7021 <= q_wait5901;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5897\ := X"0000000" & X"0";
                \$v5898\ := X"0000000" & X"1";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14407\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5897\ & "0000" & \$10734\ & "0001" & \$v5898\;
                state_var7021 <= pause_setI5899;
              end if;
            when pause_getII5912 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14405_i\ := \$$10702_brk_value\;
              \$v5910\ := \$$10698_heap_ptr_take\;
              if \$v5910\(0) = '1' then
                state_var7021 <= q_wait5909;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14405_i\;
                state_var7021 <= pause_setI5907;
              end if;
            when pause_getII5916 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14405_i\ := \$$10702_brk_value\;
              \$v5910\ := \$$10698_heap_ptr_take\;
              if \$v5910\(0) = '1' then
                state_var7021 <= q_wait5909;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14405_i\;
                state_var7021 <= pause_setI5907;
              end if;
            when pause_getII5924 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14415\ := \$$10702_brk_value\;
              \$v5922\ := \$$10702_brk_ptr_take\;
              if \$v5922\(0) = '1' then
                state_var7021 <= q_wait5921;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14415\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5919;
              end if;
            when pause_getII5929 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$10737\ := \$$10695_limit_value\;
              \$v5927\ := eclat_eq(\$10736\ & eclat_sub(\$10737\ & X"0000000" & X"1"));
              if \$v5927\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14423_forever3163312\;
              else
                \$v5926\ := \$$10702_brk_ptr_take\;
                if \$v5926\(0) = '1' then
                  state_var7021 <= q_wait5925;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5923;
                end if;
              end if;
            when pause_getII5933 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$10736\ := \$$10702_brk_value\;
              \$v5931\ := \$$10695_limit_ptr_take\;
              if \$v5931\(0) = '1' then
                state_var7021 <= q_wait5930;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5928;
              end if;
            when pause_getII5937 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$10734\ := \$$10699_symtbl_value\;
              \$v5935\ := \$$10702_brk_ptr_take\;
              if \$v5935\(0) = '1' then
                state_var7021 <= q_wait5934;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5932;
              end if;
            when pause_getII5949 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10726\ := \$$10696_ram_value\;
              \$v5945\ := \$10726\(72 to 107);
              \$v5946\ := \$v5945\(0 to 3);
              \$v5944\ := \$v5945\(4 to 35);
              case \$v5946\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14437_forever3163313\;
              when "0000" =>
                \$14445_i\ := \$v5944\(0 to 31);
                \$10731\ := \$14445_i\;
                \$v5943\ := \$$10700_pc_ptr_take\;
                if \$v5943\(0) = '1' then
                  state_var7021 <= q_wait5942;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr_write\ <= 0;
                  \$$10700_pc_write_request\ <= '1';
                  \$$10700_pc_write\ <= \$10731\;
                  state_var7021 <= pause_setI5940;
                end if;
              when others =>
                
              end case;
            when pause_getII5956 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$10721\ := \$$10696_ram_value\;
              \$v5952\ := \$10721\(0 to 35);
              \$v5953\ := \$v5952\(0 to 3);
              \$v5947\ := \$v5952\(4 to 35);
              case \$v5953\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14450_forever3163314\;
              when "0000" =>
                \$14458_i\ := \$v5947\(0 to 31);
                \$v5951\ := \$$10696_ram_ptr_take\;
                if \$v5951\(0) = '1' then
                  state_var7021 <= q_wait5950;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14458_i\));
                  state_var7021 <= pause_getI5948;
                end if;
              when others =>
                
              end case;
            when pause_getII5962 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$10720\ := \$$10698_heap_value\;
              \$v5959\ := "0000" & \$10720\;
              \$v5960\ := \$v5959\(0 to 3);
              \$v5954\ := \$v5959\(4 to 35);
              case \$v5960\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14464_forever3163315\;
              when "0000" =>
                \$14472_i\ := \$v5954\(0 to 31);
                \$v5958\ := \$$10696_ram_ptr_take\;
                if \$v5958\(0) = '1' then
                  state_var7021 <= q_wait5957;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14472_i\));
                  state_var7021 <= pause_getI5955;
                end if;
              when others =>
                
              end case;
            when pause_getII5972 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15092\ := \$$10696_ram_value\;
              \$v5969\ := \$$10696_ram_ptr_take\;
              if \$v5969\(0) = '1' then
                state_var7021 <= q_wait5968;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15090_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15076_new_rib\ & \$15091\(36 to 71) & \$15092\(72 to 107);
                state_var7021 <= pause_setI5966;
              end if;
            when pause_getII5979 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15091\ := \$$10696_ram_value\;
              \$v5975\ := "0000" & \$15070\;
              \$v5976\ := \$v5975\(0 to 3);
              \$v5970\ := \$v5975\(4 to 35);
              case \$v5976\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15106_forever3163337\;
              when "0000" =>
                \$15114_i\ := \$v5970\(0 to 31);
                \$v5974\ := \$$10696_ram_ptr_take\;
                if \$v5974\(0) = '1' then
                  state_var7021 <= q_wait5973;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$15114_i\));
                  state_var7021 <= pause_getI5971;
                end if;
              when others =>
                
              end case;
            when pause_getII5987 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$15137\ := \$$10698_heap_value\;
              \$15076_new_rib\ := "0000" & \$15137\;
              \$v5984\ := "0000" & \$15070\;
              \$v5985\ := \$v5984\(0 to 3);
              \$v5965\ := \$v5984\(4 to 35);
              case \$v5985\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15082_forever3163336\;
              when "0000" =>
                \$15090_i\ := \$v5965\(0 to 31);
                \$v5982\ := "0000" & \$15070\;
                \$v5983\ := \$v5982\(0 to 3);
                \$v5977\ := \$v5982\(4 to 35);
                case \$v5983\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$15120_forever3163338\;
                when "0000" =>
                  \$15128_i\ := \$v5977\(0 to 31);
                  \$v5981\ := \$$10696_ram_ptr_take\;
                  if \$v5981\(0) = '1' then
                    state_var7021 <= q_wait5980;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$15128_i\));
                    state_var7021 <= pause_getI5978;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII5996 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$15131\ := \$$10698_heap_value\;
              \$v5994\ := \$$10696_ram_ptr_take\;
              if \$v5994\(0) = '1' then
                state_var7021 <= q_wait5993;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5990\ := X"0000000" & X"4";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15131\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5990\ & \$15068_opnd\ & \$15071\(0 to 35);
                state_var7021 <= pause_setI5991;
              end if;
            when pause_getII6004 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15129_i\ := \$$10702_brk_value\;
              \$v6002\ := \$$10698_heap_ptr_take\;
              if \$v6002\(0) = '1' then
                state_var7021 <= q_wait6001;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$15129_i\;
                state_var7021 <= pause_setI5999;
              end if;
            when pause_getII6008 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15129_i\ := \$$10702_brk_value\;
              \$v6002\ := \$$10698_heap_ptr_take\;
              if \$v6002\(0) = '1' then
                state_var7021 <= q_wait6001;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$15129_i\;
                state_var7021 <= pause_setI5999;
              end if;
            when pause_getII6016 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15141\ := \$$10702_brk_value\;
              \$v6014\ := \$$10702_brk_ptr_take\;
              if \$v6014\(0) = '1' then
                state_var7021 <= q_wait6013;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15141\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6011;
              end if;
            when pause_getII6021 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15075\ := \$$10695_limit_value\;
              \$v6019\ := eclat_eq(\$15074\ & eclat_sub(\$15075\ & X"0000000" & X"1"));
              if \$v6019\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15149_forever3163339\;
              else
                \$v6018\ := \$$10702_brk_ptr_take\;
                if \$v6018\(0) = '1' then
                  state_var7021 <= q_wait6017;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6015;
                end if;
              end if;
            when pause_getII6025 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15074\ := \$$10702_brk_value\;
              \$v6023\ := \$$10695_limit_ptr_take\;
              if \$v6023\(0) = '1' then
                state_var7021 <= q_wait6022;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6020;
              end if;
            when pause_getII6030 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15071\ := \$$10696_ram_value\;
              \$v6027\ := \$$10702_brk_ptr_take\;
              if \$v6027\(0) = '1' then
                state_var7021 <= q_wait6026;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6024;
              end if;
            when pause_getII6036 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$15070\ := \$$10697_stack_value\;
              \$v6033\ := "0000" & \$15070\;
              \$v6034\ := \$v6033\(0 to 3);
              \$v6028\ := \$v6033\(4 to 35);
              case \$v6034\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15164_forever3163340\;
              when "0000" =>
                \$15172_i\ := \$v6028\(0 to 31);
                \$v6032\ := \$$10696_ram_ptr_take\;
                if \$v6032\(0) = '1' then
                  state_var7021 <= q_wait6031;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$15172_i\));
                  state_var7021 <= pause_getI6029;
                end if;
              when others =>
                
              end case;
            when pause_getII6047 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15063\ := \$$10696_ram_value\;
              \$v6044\ := \$15063\(36 to 71);
              \$v6045\ := \$v6044\(0 to 3);
              \$v6043\ := \$v6044\(4 to 35);
              case \$v6045\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15178_forever3163341\;
              when "0000" =>
                \$15186_i\ := \$v6043\(0 to 31);
                \$15067\ := \$15186_i\;
                \$v6042\ := \$$10697_stack_ptr_take\;
                if \$v6042\(0) = '1' then
                  state_var7021 <= q_wait6041;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$15067\;
                  state_var7021 <= pause_setI6039;
                end if;
              when others =>
                
              end case;
            when pause_getII6051 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$15062\ := \$$10697_stack_value\;
              \$v6049\ := \$$10696_ram_ptr_take\;
              if \$v6049\(0) = '1' then
                state_var7021 <= q_wait6048;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15062\));
                state_var7021 <= pause_getI6046;
              end if;
            when pause_getII6061 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14683\ := \$$10696_ram_value\;
              \$v6058\ := \$$10696_ram_ptr_take\;
              if \$v6058\(0) = '1' then
                state_var7021 <= q_wait6057;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14681_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$14667_new_rib\ & \$14682\(36 to 71) & \$14683\(72 to 107);
                state_var7021 <= pause_setI6055;
              end if;
            when pause_getII6068 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14682\ := \$$10696_ram_value\;
              \$v6064\ := "0000" & \$14661\;
              \$v6065\ := \$v6064\(0 to 3);
              \$v6059\ := \$v6064\(4 to 35);
              case \$v6065\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14697_forever3163322\;
              when "0000" =>
                \$14705_i\ := \$v6059\(0 to 31);
                \$v6063\ := \$$10696_ram_ptr_take\;
                if \$v6063\(0) = '1' then
                  state_var7021 <= q_wait6062;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14705_i\));
                  state_var7021 <= pause_getI6060;
                end if;
              when others =>
                
              end case;
            when pause_getII6076 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14728\ := \$$10698_heap_value\;
              \$14667_new_rib\ := "0000" & \$14728\;
              \$v6073\ := "0000" & \$14661\;
              \$v6074\ := \$v6073\(0 to 3);
              \$v6054\ := \$v6073\(4 to 35);
              case \$v6074\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14673_forever3163321\;
              when "0000" =>
                \$14681_i\ := \$v6054\(0 to 31);
                \$v6071\ := "0000" & \$14661\;
                \$v6072\ := \$v6071\(0 to 3);
                \$v6066\ := \$v6071\(4 to 35);
                case \$v6072\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14711_forever3163323\;
                when "0000" =>
                  \$14719_i\ := \$v6066\(0 to 31);
                  \$v6070\ := \$$10696_ram_ptr_take\;
                  if \$v6070\(0) = '1' then
                    state_var7021 <= q_wait6069;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14719_i\));
                    state_var7021 <= pause_getI6067;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII6085 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14722\ := \$$10698_heap_value\;
              \$v6083\ := \$$10696_ram_ptr_take\;
              if \$v6083\(0) = '1' then
                state_var7021 <= q_wait6082;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6079\ := X"0000000" & X"3";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14722\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v6079\ & \$14656_proc_rib\ & \$14662\(0 to 35);
                state_var7021 <= pause_setI6080;
              end if;
            when pause_getII6093 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14720_i\ := \$$10702_brk_value\;
              \$v6091\ := \$$10698_heap_ptr_take\;
              if \$v6091\(0) = '1' then
                state_var7021 <= q_wait6090;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14720_i\;
                state_var7021 <= pause_setI6088;
              end if;
            when pause_getII6097 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14720_i\ := \$$10702_brk_value\;
              \$v6091\ := \$$10698_heap_ptr_take\;
              if \$v6091\(0) = '1' then
                state_var7021 <= q_wait6090;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14720_i\;
                state_var7021 <= pause_setI6088;
              end if;
            when pause_getII6105 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14732\ := \$$10702_brk_value\;
              \$v6103\ := \$$10702_brk_ptr_take\;
              if \$v6103\(0) = '1' then
                state_var7021 <= q_wait6102;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14732\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6100;
              end if;
            when pause_getII6110 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$14666\ := \$$10695_limit_value\;
              \$v6108\ := eclat_eq(\$14665\ & eclat_sub(\$14666\ & X"0000000" & X"1"));
              if \$v6108\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14740_forever3163324\;
              else
                \$v6107\ := \$$10702_brk_ptr_take\;
                if \$v6107\(0) = '1' then
                  state_var7021 <= q_wait6106;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6104;
                end if;
              end if;
            when pause_getII6114 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14665\ := \$$10702_brk_value\;
              \$v6112\ := \$$10695_limit_ptr_take\;
              if \$v6112\(0) = '1' then
                state_var7021 <= q_wait6111;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6109;
              end if;
            when pause_getII6119 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14662\ := \$$10696_ram_value\;
              \$v6116\ := \$$10702_brk_ptr_take\;
              if \$v6116\(0) = '1' then
                state_var7021 <= q_wait6115;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6113;
              end if;
            when pause_getII6125 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$14661\ := \$$10697_stack_value\;
              \$v6122\ := "0000" & \$14661\;
              \$v6123\ := \$v6122\(0 to 3);
              \$v6117\ := \$v6122\(4 to 35);
              case \$v6123\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14755_forever3163325\;
              when "0000" =>
                \$14763_i\ := \$v6117\(0 to 31);
                \$v6121\ := \$$10696_ram_ptr_take\;
                if \$v6121\(0) = '1' then
                  state_var7021 <= q_wait6120;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14763_i\));
                  state_var7021 <= pause_getI6118;
                end if;
              when others =>
                
              end case;
            when pause_getII6133 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$14658\ := \$$10697_stack_value\;
              \$v6130\ := "0000" & \$14658\;
              \$v6131\ := \$v6130\(0 to 3);
              \$v6129\ := \$v6130\(4 to 35);
              case \$v6131\ is
              when "0001" =>
                \$14659\ := eclat_false;
              when "0000" =>
                \$14766_i\ := \$v6129\(0 to 31);
                \$14659\ := eclat_if(eclat_ge(\$14766_i\ & X"0000000" & X"0") & eclat_lt(\$14766_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v6128\ := \$14659\;
              if \$v6128\(0) = '1' then
                \$v6127\ := \$$10697_stack_ptr_take\;
                if \$v6127\(0) = '1' then
                  state_var7021 <= q_wait6126;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI6124;
                end if;
              else
                \$14511_loop311_result\ := eclat_unit;
                \$14481_decode_loop310_result\ := \$14511_loop311_result\;
                \$v5964\ := \$$10698_heap_ptr_take\;
                if \$v5964\(0) = '1' then
                  state_var7021 <= q_wait5963;
                else
                  \$$10698_heap_ptr_take\(0) := '1';
                  \$$10698_heap_ptr\ <= 0;
                  state_var7021 <= pause_getI5961;
                end if;
              end if;
            when pause_getII6137 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14772\ := \$$10698_heap_value\;
              \$14656_proc_rib\ := "0000" & \$14772\;
              \$v6135\ := \$$10697_stack_ptr_take\;
              if \$v6135\(0) = '1' then
                state_var7021 <= q_wait6134;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6132;
              end if;
            when pause_getII6147 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14770\ := \$$10698_heap_value\;
              \$v6145\ := \$$10696_ram_ptr_take\;
              if \$v6145\(0) = '1' then
                state_var7021 <= q_wait6144;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6140\ := X"0000000" & X"0";
                \$v6141\ := X"0000000" & X"1";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14770\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$14652_code_proc_rib\ & "0000" & \$v6140\ & "0001" & \$v6141\;
                state_var7021 <= pause_setI6142;
              end if;
            when pause_getII6155 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14768_i\ := \$$10702_brk_value\;
              \$v6153\ := \$$10698_heap_ptr_take\;
              if \$v6153\(0) = '1' then
                state_var7021 <= q_wait6152;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14768_i\;
                state_var7021 <= pause_setI6150;
              end if;
            when pause_getII6159 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14768_i\ := \$$10702_brk_value\;
              \$v6153\ := \$$10698_heap_ptr_take\;
              if \$v6153\(0) = '1' then
                state_var7021 <= q_wait6152;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14768_i\;
                state_var7021 <= pause_setI6150;
              end if;
            when pause_getII6167 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14777\ := \$$10702_brk_value\;
              \$v6165\ := \$$10702_brk_ptr_take\;
              if \$v6165\(0) = '1' then
                state_var7021 <= q_wait6164;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14777\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6162;
              end if;
            when pause_getII6172 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$14655\ := \$$10695_limit_value\;
              \$v6170\ := eclat_eq(\$14654\ & eclat_sub(\$14655\ & X"0000000" & X"1"));
              if \$v6170\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14785_forever3163326\;
              else
                \$v6169\ := \$$10702_brk_ptr_take\;
                if \$v6169\(0) = '1' then
                  state_var7021 <= q_wait6168;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6166;
                end if;
              end if;
            when pause_getII6176 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14654\ := \$$10702_brk_value\;
              \$v6174\ := \$$10695_limit_ptr_take\;
              if \$v6174\(0) = '1' then
                state_var7021 <= q_wait6173;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6171;
              end if;
            when pause_getII6180 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14799\ := \$$10698_heap_value\;
              \$14652_code_proc_rib\ := "0000" & \$14799\;
              \$v6178\ := \$$10702_brk_ptr_take\;
              if \$v6178\(0) = '1' then
                state_var7021 <= q_wait6177;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6175;
              end if;
            when pause_getII6189 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14797\ := \$$10698_heap_value\;
              \$v6187\ := \$$10696_ram_ptr_take\;
              if \$v6187\(0) = '1' then
                state_var7021 <= q_wait6186;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6183\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14797\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$14533_opnd\ & "0001" & \$v6183\ & \$14648_ty\;
                state_var7021 <= pause_setI6184;
              end if;
            when pause_getII6197 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14795_i\ := \$$10702_brk_value\;
              \$v6195\ := \$$10698_heap_ptr_take\;
              if \$v6195\(0) = '1' then
                state_var7021 <= q_wait6194;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14795_i\;
                state_var7021 <= pause_setI6192;
              end if;
            when pause_getII6201 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14795_i\ := \$$10702_brk_value\;
              \$v6195\ := \$$10698_heap_ptr_take\;
              if \$v6195\(0) = '1' then
                state_var7021 <= q_wait6194;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14795_i\;
                state_var7021 <= pause_setI6192;
              end if;
            when pause_getII6209 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14803\ := \$$10702_brk_value\;
              \$v6207\ := \$$10702_brk_ptr_take\;
              if \$v6207\(0) = '1' then
                state_var7021 <= q_wait6206;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14803\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6204;
              end if;
            when pause_getII6214 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$14651\ := \$$10695_limit_value\;
              \$v6212\ := eclat_eq(\$14650\ & eclat_sub(\$14651\ & X"0000000" & X"1"));
              if \$v6212\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14811_forever3163327\;
              else
                \$v6211\ := \$$10702_brk_ptr_take\;
                if \$v6211\(0) = '1' then
                  state_var7021 <= q_wait6210;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6208;
                end if;
              end if;
            when pause_getII6218 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14650\ := \$$10702_brk_value\;
              \$v6216\ := \$$10695_limit_ptr_take\;
              if \$v6216\(0) = '1' then
                state_var7021 <= q_wait6215;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6213;
              end if;
            when pause_getII6229 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14643\ := \$$10696_ram_value\;
              \$v6226\ := \$14643\(36 to 71);
              \$v6227\ := \$v6226\(0 to 3);
              \$v6225\ := \$v6226\(4 to 35);
              case \$v6227\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14826_forever3163328\;
              when "0000" =>
                \$14834_i\ := \$v6225\(0 to 31);
                \$14647\ := \$14834_i\;
                \$v6224\ := \$$10697_stack_ptr_take\;
                if \$v6224\(0) = '1' then
                  state_var7021 <= q_wait6223;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$14647\;
                  state_var7021 <= pause_setI6221;
                end if;
              when others =>
                
              end case;
            when pause_getII6233 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$14642\ := \$$10697_stack_value\;
              \$v6231\ := \$$10696_ram_ptr_take\;
              if \$v6231\(0) = '1' then
                state_var7021 <= q_wait6230;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14642\));
                state_var7021 <= pause_getI6228;
              end if;
            when pause_getII6243 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14558\ := \$$10696_ram_value\;
              \$v6240\ := \$$10696_ram_ptr_take\;
              if \$v6240\(0) = '1' then
                state_var7021 <= q_wait6239;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14556_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$14542_new_rib\ & \$14557\(36 to 71) & \$14558\(72 to 107);
                state_var7021 <= pause_setI6237;
              end if;
            when pause_getII6250 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14557\ := \$$10696_ram_value\;
              \$v6246\ := "0000" & \$14536\;
              \$v6247\ := \$v6246\(0 to 3);
              \$v6241\ := \$v6246\(4 to 35);
              case \$v6247\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14572_forever3163317\;
              when "0000" =>
                \$14580_i\ := \$v6241\(0 to 31);
                \$v6245\ := \$$10696_ram_ptr_take\;
                if \$v6245\(0) = '1' then
                  state_var7021 <= q_wait6244;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14580_i\));
                  state_var7021 <= pause_getI6242;
                end if;
              when others =>
                
              end case;
            when pause_getII6258 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14603\ := \$$10698_heap_value\;
              \$14542_new_rib\ := "0000" & \$14603\;
              \$v6255\ := "0000" & \$14536\;
              \$v6256\ := \$v6255\(0 to 3);
              \$v6236\ := \$v6255\(4 to 35);
              case \$v6256\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14548_forever3163316\;
              when "0000" =>
                \$14556_i\ := \$v6236\(0 to 31);
                \$v6253\ := "0000" & \$14536\;
                \$v6254\ := \$v6253\(0 to 3);
                \$v6248\ := \$v6253\(4 to 35);
                case \$v6254\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$14586_forever3163318\;
                when "0000" =>
                  \$14594_i\ := \$v6248\(0 to 31);
                  \$v6252\ := \$$10696_ram_ptr_take\;
                  if \$v6252\(0) = '1' then
                    state_var7021 <= q_wait6251;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$14594_i\));
                    state_var7021 <= pause_getI6249;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_getII6267 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$14597\ := \$$10698_heap_value\;
              \$v6265\ := \$$10696_ram_ptr_take\;
              if \$v6265\(0) = '1' then
                state_var7021 <= q_wait6264;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6261\ := eclat_if(eclat_lt(X"0000000" & X"0" & \$14511_loop311_arg\(0 to 31)) & eclat_sub(\$14511_loop311_arg\(0 to 31) & X"0000000" & X"1") & X"0000000" & X"0");
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14597\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v6261\ & \$14533_opnd\ & \$14537\(0 to 35);
                state_var7021 <= pause_setI6262;
              end if;
            when pause_getII6275 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14595_i\ := \$$10702_brk_value\;
              \$v6273\ := \$$10698_heap_ptr_take\;
              if \$v6273\(0) = '1' then
                state_var7021 <= q_wait6272;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14595_i\;
                state_var7021 <= pause_setI6270;
              end if;
            when pause_getII6279 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14595_i\ := \$$10702_brk_value\;
              \$v6273\ := \$$10698_heap_ptr_take\;
              if \$v6273\(0) = '1' then
                state_var7021 <= q_wait6272;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14595_i\;
                state_var7021 <= pause_setI6270;
              end if;
            when pause_getII6287 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14609\ := \$$10702_brk_value\;
              \$v6285\ := \$$10702_brk_ptr_take\;
              if \$v6285\(0) = '1' then
                state_var7021 <= q_wait6284;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14609\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6282;
              end if;
            when pause_getII6292 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$14541\ := \$$10695_limit_value\;
              \$v6290\ := eclat_eq(\$14540\ & eclat_sub(\$14541\ & X"0000000" & X"1"));
              if \$v6290\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14617_forever3163319\;
              else
                \$v6289\ := \$$10702_brk_ptr_take\;
                if \$v6289\(0) = '1' then
                  state_var7021 <= q_wait6288;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6286;
                end if;
              end if;
            when pause_getII6296 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$14540\ := \$$10702_brk_value\;
              \$v6294\ := \$$10695_limit_ptr_take\;
              if \$v6294\(0) = '1' then
                state_var7021 <= q_wait6293;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6291;
              end if;
            when pause_getII6301 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14537\ := \$$10696_ram_value\;
              \$v6298\ := \$$10702_brk_ptr_take\;
              if \$v6298\(0) = '1' then
                state_var7021 <= q_wait6297;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6295;
              end if;
            when pause_getII6307 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$14536\ := \$$10697_stack_value\;
              \$v6304\ := "0000" & \$14536\;
              \$v6305\ := \$v6304\(0 to 3);
              \$v6299\ := \$v6304\(4 to 35);
              case \$v6305\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$14632_forever3163320\;
              when "0000" =>
                \$14640_i\ := \$v6299\(0 to 31);
                \$v6303\ := \$$10696_ram_ptr_take\;
                if \$v6303\(0) = '1' then
                  state_var7021 <= q_wait6302;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$14640_i\));
                  state_var7021 <= pause_getI6300;
                end if;
              when others =>
                
              end case;
            when pause_getII6313 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14974\ := \$$10696_ram_value\;
              \$14533_opnd\ := \$14974\(0 to 35);
              \$v6310\ := eclat_lt(X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31));
              if \$v6310\(0) = '1' then
                \$v6235\ := \$$10697_stack_ptr_take\;
                if \$v6235\(0) = '1' then
                  state_var7021 <= q_wait6234;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI6232;
                end if;
              else
                \$v6309\ := \$$10697_stack_ptr_take\;
                if \$v6309\(0) = '1' then
                  state_var7021 <= q_wait6308;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI6306;
                end if;
              end if;
            when pause_getII6320 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15005\ := \$$10696_ram_value\;
              \$14996_list_tail2653334_arg\ := \$15005\(36 to 71) & eclat_sub(\$14996_list_tail2653334_arg\(36 to 67) & X"0000000" & X"1") & eclat_unit;
              state_var7021 <= \$14996_list_tail2653334\;
            when pause_getII6327 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$14972\ := \$$10699_symtbl_value\;
              \$14996_list_tail2653334_arg\ := "0000" & \$14972\ & \$14511_loop311_arg\(32 to 63) & eclat_unit;
              state_var7021 <= \$14996_list_tail2653334\;
            when pause_getII6338 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14948\ := \$$10701_pos_value\;
              \$v6336\ := \$$10701_pos_ptr_take\;
              if \$v6336\(0) = '1' then
                state_var7021 <= q_wait6335;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$14948\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6333;
              end if;
            when pause_getII6342 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14947\ := \$$10701_pos_value\;
              \$v6340\ := \$$10701_pos_ptr_take\;
              if \$v6340\(0) = '1' then
                state_var7021 <= q_wait6339;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6337;
              end if;
            when pause_getII6347 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14841\ := \$$10696_ram_value\;
              \$14533_opnd\ := \$14841\(0 to 35);
              \$v6310\ := eclat_lt(X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31));
              if \$v6310\(0) = '1' then
                \$v6235\ := \$$10697_stack_ptr_take\;
                if \$v6235\(0) = '1' then
                  state_var7021 <= q_wait6234;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI6232;
                end if;
              else
                \$v6309\ := \$$10697_stack_ptr_take\;
                if \$v6309\(0) = '1' then
                  state_var7021 <= q_wait6308;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI6306;
                end if;
              end if;
            when pause_getII6354 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$14872\ := \$$10696_ram_value\;
              \$14863_list_tail2653331_arg\ := \$14872\(36 to 71) & eclat_sub(\$14863_list_tail2653331_arg\(36 to 67) & X"0000000" & X"1") & eclat_unit;
              state_var7021 <= \$14863_list_tail2653331\;
            when pause_getII6361 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$14839\ := \$$10699_symtbl_value\;
              \$14863_list_tail2653331_arg\ := "0000" & \$14839\ & \$14837\ & eclat_unit;
              state_var7021 <= \$14863_list_tail2653331\;
            when pause_getII6370 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14912\ := \$$10701_pos_value\;
              \$v6368\ := \$$10701_pos_ptr_take\;
              if \$v6368\(0) = '1' then
                state_var7021 <= q_wait6367;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$14912\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6365;
              end if;
            when pause_getII6374 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14911\ := \$$10701_pos_value\;
              \$v6372\ := \$$10701_pos_ptr_take\;
              if \$v6372\(0) = '1' then
                state_var7021 <= q_wait6371;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6369;
              end if;
            when pause_getII6386 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$15037\ := \$$10697_stack_value\;
              \$v6384\ := \$$10696_ram_ptr_take\;
              if \$v6384\(0) = '1' then
                state_var7021 <= q_wait6383;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6379\ := \$14511_loop311_arg\(0 to 31);
                \$v6380\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15037\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v6379\ & "0000" & \$15035\ & "0001" & \$v6380\;
                state_var7021 <= pause_setI6381;
              end if;
            when pause_getII6394 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$15035\ := \$$10697_stack_value\;
              \$v6392\ := \$$10697_stack_ptr_take\;
              if \$v6392\(0) = '1' then
                state_var7021 <= q_wait6391;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$15034_i\;
                state_var7021 <= pause_setI6389;
              end if;
            when pause_getII6398 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15034_i\ := \$$10702_brk_value\;
              \$v6396\ := \$$10697_stack_ptr_take\;
              if \$v6396\(0) = '1' then
                state_var7021 <= q_wait6395;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6393;
              end if;
            when pause_getII6402 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15034_i\ := \$$10702_brk_value\;
              \$v6396\ := \$$10697_stack_ptr_take\;
              if \$v6396\(0) = '1' then
                state_var7021 <= q_wait6395;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6393;
              end if;
            when pause_getII6410 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15043\ := \$$10702_brk_value\;
              \$v6408\ := \$$10702_brk_ptr_take\;
              if \$v6408\(0) = '1' then
                state_var7021 <= q_wait6407;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15043\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6405;
              end if;
            when pause_getII6415 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15033\ := \$$10695_limit_value\;
              \$v6413\ := eclat_eq(\$15032\ & eclat_sub(\$15033\ & X"0000000" & X"1"));
              if \$v6413\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15051_forever3163335\;
              else
                \$v6412\ := \$$10702_brk_ptr_take\;
                if \$v6412\(0) = '1' then
                  state_var7021 <= q_wait6411;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6409;
                end if;
              end if;
            when pause_getII6419 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15032\ := \$$10702_brk_value\;
              \$v6417\ := \$$10695_limit_ptr_take\;
              if \$v6417\(0) = '1' then
                state_var7021 <= q_wait6416;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6414;
              end if;
            when pause_getII6430 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14499\ := \$$10701_pos_value\;
              \$v6428\ := \$$10701_pos_ptr_take\;
              if \$v6428\(0) = '1' then
                state_var7021 <= q_wait6427;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$14499\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6425;
              end if;
            when pause_getII6434 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14498\ := \$$10701_pos_value\;
              \$v6432\ := \$$10701_pos_ptr_take\;
              if \$v6432\(0) = '1' then
                state_var7021 <= q_wait6431;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6429;
              end if;
            when pause_getII6438 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15650\ := \$$10699_symtbl_value\;
              \$15217_loop1312_arg\ := eclat_sub(\$15217_loop1312_arg\(0 to 31) & X"0000000" & X"1") & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var7021 <= \$15217_loop1312\;
            when pause_getII6447 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15648\ := \$$10699_symtbl_value\;
              \$v6445\ := \$$10696_ram_ptr_take\;
              if \$v6445\(0) = '1' then
                state_var7021 <= q_wait6444;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6441\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15648\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15642_end_rib\ & "0000" & \$15621\ & "0001" & \$v6441\;
                state_var7021 <= pause_setI6442;
              end if;
            when pause_getII6455 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15646_i\ := \$$10702_brk_value\;
              \$v6453\ := \$$10699_symtbl_ptr_take\;
              if \$v6453\(0) = '1' then
                state_var7021 <= q_wait6452;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15646_i\;
                state_var7021 <= pause_setI6450;
              end if;
            when pause_getII6459 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15646_i\ := \$$10702_brk_value\;
              \$v6453\ := \$$10699_symtbl_ptr_take\;
              if \$v6453\(0) = '1' then
                state_var7021 <= q_wait6452;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15646_i\;
                state_var7021 <= pause_setI6450;
              end if;
            when pause_getII6467 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15655\ := \$$10702_brk_value\;
              \$v6465\ := \$$10702_brk_ptr_take\;
              if \$v6465\(0) = '1' then
                state_var7021 <= q_wait6464;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15655\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6462;
              end if;
            when pause_getII6472 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15645\ := \$$10695_limit_value\;
              \$v6470\ := eclat_eq(\$15644\ & eclat_sub(\$15645\ & X"0000000" & X"1"));
              if \$v6470\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15663_forever3163356\;
              else
                \$v6469\ := \$$10702_brk_ptr_take\;
                if \$v6469\(0) = '1' then
                  state_var7021 <= q_wait6468;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6466;
                end if;
              end if;
            when pause_getII6476 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15644\ := \$$10702_brk_value\;
              \$v6474\ := \$$10695_limit_ptr_take\;
              if \$v6474\(0) = '1' then
                state_var7021 <= q_wait6473;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6471;
              end if;
            when pause_getII6480 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15673\ := \$$10699_symtbl_value\;
              \$15642_end_rib\ := "0000" & \$15673\;
              \$v6478\ := \$$10702_brk_ptr_take\;
              if \$v6478\(0) = '1' then
                state_var7021 <= q_wait6477;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6475;
              end if;
            when pause_getII6490 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15640\ := \$$10699_symtbl_value\;
              \$v6488\ := \$$10696_ram_ptr_take\;
              if \$v6488\(0) = '1' then
                state_var7021 <= q_wait6487;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6483\ := X"0000000" & X"2";
                \$v6484\ := X"0000000" & X"2";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15640\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v6483\ & \$15634_str_rib\ & "0001" & \$v6484\;
                state_var7021 <= pause_setI6485;
              end if;
            when pause_getII6498 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15638_i\ := \$$10702_brk_value\;
              \$v6496\ := \$$10699_symtbl_ptr_take\;
              if \$v6496\(0) = '1' then
                state_var7021 <= q_wait6495;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15638_i\;
                state_var7021 <= pause_setI6493;
              end if;
            when pause_getII6502 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15638_i\ := \$$10702_brk_value\;
              \$v6496\ := \$$10699_symtbl_ptr_take\;
              if \$v6496\(0) = '1' then
                state_var7021 <= q_wait6495;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15638_i\;
                state_var7021 <= pause_setI6493;
              end if;
            when pause_getII6510 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15678\ := \$$10702_brk_value\;
              \$v6508\ := \$$10702_brk_ptr_take\;
              if \$v6508\(0) = '1' then
                state_var7021 <= q_wait6507;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15678\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6505;
              end if;
            when pause_getII6515 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15637\ := \$$10695_limit_value\;
              \$v6513\ := eclat_eq(\$15636\ & eclat_sub(\$15637\ & X"0000000" & X"1"));
              if \$v6513\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15686_forever3163357\;
              else
                \$v6512\ := \$$10702_brk_ptr_take\;
                if \$v6512\(0) = '1' then
                  state_var7021 <= q_wait6511;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6509;
                end if;
              end if;
            when pause_getII6519 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15636\ := \$$10702_brk_value\;
              \$v6517\ := \$$10695_limit_ptr_take\;
              if \$v6517\(0) = '1' then
                state_var7021 <= q_wait6516;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6514;
              end if;
            when pause_getII6523 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15696\ := \$$10699_symtbl_value\;
              \$15634_str_rib\ := "0000" & \$15696\;
              \$v6521\ := \$$10702_brk_ptr_take\;
              if \$v6521\(0) = '1' then
                state_var7021 <= q_wait6520;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6518;
              end if;
            when pause_getII6533 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15632\ := \$$10699_symtbl_value\;
              \$v6531\ := \$$10696_ram_ptr_take\;
              if \$v6531\(0) = '1' then
                state_var7021 <= q_wait6530;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6526\ := X"0000000" & X"0";
                \$v6527\ := X"0000000" & X"3";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15632\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v6526\ & "0001" & \$15622\ & "0001" & \$v6527\;
                state_var7021 <= pause_setI6528;
              end if;
            when pause_getII6541 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15630_i\ := \$$10702_brk_value\;
              \$v6539\ := \$$10699_symtbl_ptr_take\;
              if \$v6539\(0) = '1' then
                state_var7021 <= q_wait6538;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15630_i\;
                state_var7021 <= pause_setI6536;
              end if;
            when pause_getII6545 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15630_i\ := \$$10702_brk_value\;
              \$v6539\ := \$$10699_symtbl_ptr_take\;
              if \$v6539\(0) = '1' then
                state_var7021 <= q_wait6538;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15630_i\;
                state_var7021 <= pause_setI6536;
              end if;
            when pause_getII6553 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15702\ := \$$10702_brk_value\;
              \$v6551\ := \$$10702_brk_ptr_take\;
              if \$v6551\(0) = '1' then
                state_var7021 <= q_wait6550;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15702\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6548;
              end if;
            when pause_getII6558 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15629\ := \$$10695_limit_value\;
              \$v6556\ := eclat_eq(\$15628\ & eclat_sub(\$15629\ & X"0000000" & X"1"));
              if \$v6556\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15710_forever3163358\;
              else
                \$v6555\ := \$$10702_brk_ptr_take\;
                if \$v6555\(0) = '1' then
                  state_var7021 <= q_wait6554;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6552;
                end if;
              end if;
            when pause_getII6562 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15628\ := \$$10702_brk_value\;
              \$v6560\ := \$$10695_limit_ptr_take\;
              if \$v6560\(0) = '1' then
                state_var7021 <= q_wait6559;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6557;
              end if;
            when pause_getII6567 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15734\ := \$$10696_ram_value\;
              \$15724_len_aux3143361_arg\ := \$15734\(36 to 71) & eclat_add(\$15724_len_aux3143361_arg\(36 to 67) & X"0000000" & X"1") & eclat_unit;
              state_var7021 <= \$15724_len_aux3143361\;
            when pause_getII6586 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15755\ := \$$10696_ram_value\;
              \$v6582\ := \$15755\(72 to 107);
              \$v6583\ := \$v6582\(0 to 3);
              \$v6573\ := \$v6582\(4 to 35);
              case \$v6583\ is
              when "0001" =>
                \$15760_i\ := \$v6573\(0 to 31);
                \$v6577\ := X"0000000" & X"0";
                \$v6575\ := "0001" & \$v6577\;
                \$v6576\ := \$v6575\(0 to 3);
                \$v6574\ := \$v6575\(4 to 35);
                case \$v6576\ is
                when "0000" =>
                  \$15733\ := eclat_false;
                when "0001" =>
                  \$15763_j\ := \$v6574\(0 to 31);
                  \$15733\ := eclat_eq(\$15760_i\ & \$15763_j\);
                when others =>
                  
                end case;
                \$v6572\ := \$15733\;
                if \$v6572\(0) = '1' then
                  \$v6570\ := \$15724_len_aux3143361_arg\(0 to 35);
                  \$v6571\ := \$v6570\(0 to 3);
                  \$v6565\ := \$v6570\(4 to 35);
                  case \$v6571\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15746_forever3163359\;
                  when "0000" =>
                    \$15754_i\ := \$v6565\(0 to 31);
                    \$v6569\ := \$$10696_ram_ptr_take\;
                    if \$v6569\(0) = '1' then
                      state_var7021 <= q_wait6568;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15754_i\));
                      state_var7021 <= pause_getI6566;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15724_len_aux3143361_result\ := \$15724_len_aux3143361_arg\(36 to 67);
                  \$15622\ := \$15724_len_aux3143361_result\;
                  \$v6564\ := \$$10702_brk_ptr_take\;
                  if \$v6564\(0) = '1' then
                    state_var7021 <= q_wait6563;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6561;
                  end if;
                end if;
              when "0000" =>
                \$15764_i\ := \$v6573\(0 to 31);
                \$v6581\ := X"0000000" & X"0";
                \$v6579\ := "0001" & \$v6581\;
                \$v6580\ := \$v6579\(0 to 3);
                \$v6578\ := \$v6579\(4 to 35);
                case \$v6580\ is
                when "0001" =>
                  \$15733\ := eclat_false;
                when "0000" =>
                  \$15767_j\ := \$v6578\(0 to 31);
                  \$15733\ := eclat_eq(\$15764_i\ & \$15767_j\);
                when others =>
                  
                end case;
                \$v6572\ := \$15733\;
                if \$v6572\(0) = '1' then
                  \$v6570\ := \$15724_len_aux3143361_arg\(0 to 35);
                  \$v6571\ := \$v6570\(0 to 3);
                  \$v6565\ := \$v6570\(4 to 35);
                  case \$v6571\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15746_forever3163359\;
                  when "0000" =>
                    \$15754_i\ := \$v6565\(0 to 31);
                    \$v6569\ := \$$10696_ram_ptr_take\;
                    if \$v6569\(0) = '1' then
                      state_var7021 <= q_wait6568;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15754_i\));
                      state_var7021 <= pause_getI6566;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15724_len_aux3143361_result\ := \$15724_len_aux3143361_arg\(36 to 67);
                  \$15622\ := \$15724_len_aux3143361_result\;
                  \$v6564\ := \$$10702_brk_ptr_take\;
                  if \$v6564\(0) = '1' then
                    state_var7021 <= q_wait6563;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6561;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII6597 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15621\ := \$$10699_symtbl_value\;
              \$v6595\ := X"0000000" & X"0";
              \$15724_len_aux3143361_arg\ := "0000" & \$v6595\ & X"0000000" & X"0" & eclat_unit;
              state_var7021 <= \$15724_len_aux3143361\;
            when pause_getII6602 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15483\ := \$$10699_symtbl_value\;
              \$v6600\ := X"0000000" & X"0";
              \$15240_loop23133355_arg\ := "0000" & \$v6600\ & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var7021 <= \$15240_loop23133355\;
            when pause_getII6611 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15481\ := \$$10699_symtbl_value\;
              \$v6609\ := \$$10696_ram_ptr_take\;
              if \$v6609\(0) = '1' then
                state_var7021 <= q_wait6608;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6605\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15481\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15475_end_rib\ & "0000" & \$15454\ & "0001" & \$v6605\;
                state_var7021 <= pause_setI6606;
              end if;
            when pause_getII6619 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15479_i\ := \$$10702_brk_value\;
              \$v6617\ := \$$10699_symtbl_ptr_take\;
              if \$v6617\(0) = '1' then
                state_var7021 <= q_wait6616;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15479_i\;
                state_var7021 <= pause_setI6614;
              end if;
            when pause_getII6623 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15479_i\ := \$$10702_brk_value\;
              \$v6617\ := \$$10699_symtbl_ptr_take\;
              if \$v6617\(0) = '1' then
                state_var7021 <= q_wait6616;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15479_i\;
                state_var7021 <= pause_setI6614;
              end if;
            when pause_getII6631 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15488\ := \$$10702_brk_value\;
              \$v6629\ := \$$10702_brk_ptr_take\;
              if \$v6629\(0) = '1' then
                state_var7021 <= q_wait6628;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15488\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6626;
              end if;
            when pause_getII6636 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15478\ := \$$10695_limit_value\;
              \$v6634\ := eclat_eq(\$15477\ & eclat_sub(\$15478\ & X"0000000" & X"1"));
              if \$v6634\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15496_forever3163349\;
              else
                \$v6633\ := \$$10702_brk_ptr_take\;
                if \$v6633\(0) = '1' then
                  state_var7021 <= q_wait6632;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6630;
                end if;
              end if;
            when pause_getII6640 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15477\ := \$$10702_brk_value\;
              \$v6638\ := \$$10695_limit_ptr_take\;
              if \$v6638\(0) = '1' then
                state_var7021 <= q_wait6637;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6635;
              end if;
            when pause_getII6644 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15506\ := \$$10699_symtbl_value\;
              \$15475_end_rib\ := "0000" & \$15506\;
              \$v6642\ := \$$10702_brk_ptr_take\;
              if \$v6642\(0) = '1' then
                state_var7021 <= q_wait6641;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6639;
              end if;
            when pause_getII6654 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15473\ := \$$10699_symtbl_value\;
              \$v6652\ := \$$10696_ram_ptr_take\;
              if \$v6652\(0) = '1' then
                state_var7021 <= q_wait6651;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6647\ := X"0000000" & X"2";
                \$v6648\ := X"0000000" & X"2";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15473\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v6647\ & \$15467_str_rib\ & "0001" & \$v6648\;
                state_var7021 <= pause_setI6649;
              end if;
            when pause_getII6662 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15471_i\ := \$$10702_brk_value\;
              \$v6660\ := \$$10699_symtbl_ptr_take\;
              if \$v6660\(0) = '1' then
                state_var7021 <= q_wait6659;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15471_i\;
                state_var7021 <= pause_setI6657;
              end if;
            when pause_getII6666 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15471_i\ := \$$10702_brk_value\;
              \$v6660\ := \$$10699_symtbl_ptr_take\;
              if \$v6660\(0) = '1' then
                state_var7021 <= q_wait6659;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15471_i\;
                state_var7021 <= pause_setI6657;
              end if;
            when pause_getII6674 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15511\ := \$$10702_brk_value\;
              \$v6672\ := \$$10702_brk_ptr_take\;
              if \$v6672\(0) = '1' then
                state_var7021 <= q_wait6671;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15511\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6669;
              end if;
            when pause_getII6679 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15470\ := \$$10695_limit_value\;
              \$v6677\ := eclat_eq(\$15469\ & eclat_sub(\$15470\ & X"0000000" & X"1"));
              if \$v6677\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15519_forever3163350\;
              else
                \$v6676\ := \$$10702_brk_ptr_take\;
                if \$v6676\(0) = '1' then
                  state_var7021 <= q_wait6675;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6673;
                end if;
              end if;
            when pause_getII6683 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15469\ := \$$10702_brk_value\;
              \$v6681\ := \$$10695_limit_ptr_take\;
              if \$v6681\(0) = '1' then
                state_var7021 <= q_wait6680;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6678;
              end if;
            when pause_getII6687 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15529\ := \$$10699_symtbl_value\;
              \$15467_str_rib\ := "0000" & \$15529\;
              \$v6685\ := \$$10702_brk_ptr_take\;
              if \$v6685\(0) = '1' then
                state_var7021 <= q_wait6684;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6682;
              end if;
            when pause_getII6696 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15465\ := \$$10699_symtbl_value\;
              \$v6694\ := \$$10696_ram_ptr_take\;
              if \$v6694\(0) = '1' then
                state_var7021 <= q_wait6693;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6690\ := X"0000000" & X"3";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15465\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15240_loop23133355_arg\(0 to 35) & "0001" & \$15455\ & "0001" & \$v6690\;
                state_var7021 <= pause_setI6691;
              end if;
            when pause_getII6704 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15463_i\ := \$$10702_brk_value\;
              \$v6702\ := \$$10699_symtbl_ptr_take\;
              if \$v6702\(0) = '1' then
                state_var7021 <= q_wait6701;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15463_i\;
                state_var7021 <= pause_setI6699;
              end if;
            when pause_getII6708 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15463_i\ := \$$10702_brk_value\;
              \$v6702\ := \$$10699_symtbl_ptr_take\;
              if \$v6702\(0) = '1' then
                state_var7021 <= q_wait6701;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15463_i\;
                state_var7021 <= pause_setI6699;
              end if;
            when pause_getII6716 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15534\ := \$$10702_brk_value\;
              \$v6714\ := \$$10702_brk_ptr_take\;
              if \$v6714\(0) = '1' then
                state_var7021 <= q_wait6713;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15534\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6711;
              end if;
            when pause_getII6721 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15462\ := \$$10695_limit_value\;
              \$v6719\ := eclat_eq(\$15457\ & eclat_sub(\$15462\ & X"0000000" & X"1"));
              if \$v6719\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15542_forever3163351\;
              else
                \$v6718\ := \$$10702_brk_ptr_take\;
                if \$v6718\(0) = '1' then
                  state_var7021 <= q_wait6717;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6715;
                end if;
              end if;
            when pause_getII6725 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15457\ := \$$10702_brk_value\;
              \$v6723\ := \$$10695_limit_ptr_take\;
              if \$v6723\(0) = '1' then
                state_var7021 <= q_wait6722;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6720;
              end if;
            when pause_getII6730 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15565\ := \$$10696_ram_value\;
              \$15555_len_aux3143354_arg\ := \$15565\(36 to 71) & eclat_add(\$15555_len_aux3143354_arg\(36 to 67) & X"0000000" & X"1") & eclat_unit;
              state_var7021 <= \$15555_len_aux3143354\;
            when pause_getII6749 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15586\ := \$$10696_ram_value\;
              \$v6745\ := \$15586\(72 to 107);
              \$v6746\ := \$v6745\(0 to 3);
              \$v6736\ := \$v6745\(4 to 35);
              case \$v6746\ is
              when "0001" =>
                \$15591_i\ := \$v6736\(0 to 31);
                \$v6740\ := X"0000000" & X"0";
                \$v6738\ := "0001" & \$v6740\;
                \$v6739\ := \$v6738\(0 to 3);
                \$v6737\ := \$v6738\(4 to 35);
                case \$v6739\ is
                when "0000" =>
                  \$15564\ := eclat_false;
                when "0001" =>
                  \$15594_j\ := \$v6737\(0 to 31);
                  \$15564\ := eclat_eq(\$15591_i\ & \$15594_j\);
                when others =>
                  
                end case;
                \$v6735\ := \$15564\;
                if \$v6735\(0) = '1' then
                  \$v6733\ := \$15555_len_aux3143354_arg\(0 to 35);
                  \$v6734\ := \$v6733\(0 to 3);
                  \$v6728\ := \$v6733\(4 to 35);
                  case \$v6734\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15577_forever3163352\;
                  when "0000" =>
                    \$15585_i\ := \$v6728\(0 to 31);
                    \$v6732\ := \$$10696_ram_ptr_take\;
                    if \$v6732\(0) = '1' then
                      state_var7021 <= q_wait6731;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15585_i\));
                      state_var7021 <= pause_getI6729;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15555_len_aux3143354_result\ := \$15555_len_aux3143354_arg\(36 to 67);
                  \$15455\ := \$15555_len_aux3143354_result\;
                  \$v6727\ := \$$10702_brk_ptr_take\;
                  if \$v6727\(0) = '1' then
                    state_var7021 <= q_wait6726;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6724;
                  end if;
                end if;
              when "0000" =>
                \$15595_i\ := \$v6736\(0 to 31);
                \$v6744\ := X"0000000" & X"0";
                \$v6742\ := "0001" & \$v6744\;
                \$v6743\ := \$v6742\(0 to 3);
                \$v6741\ := \$v6742\(4 to 35);
                case \$v6743\ is
                when "0001" =>
                  \$15564\ := eclat_false;
                when "0000" =>
                  \$15598_j\ := \$v6741\(0 to 31);
                  \$15564\ := eclat_eq(\$15595_i\ & \$15598_j\);
                when others =>
                  
                end case;
                \$v6735\ := \$15564\;
                if \$v6735\(0) = '1' then
                  \$v6733\ := \$15555_len_aux3143354_arg\(0 to 35);
                  \$v6734\ := \$v6733\(0 to 3);
                  \$v6728\ := \$v6733\(4 to 35);
                  case \$v6734\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15577_forever3163352\;
                  when "0000" =>
                    \$15585_i\ := \$v6728\(0 to 31);
                    \$v6732\ := \$$10696_ram_ptr_take\;
                    if \$v6732\(0) = '1' then
                      state_var7021 <= q_wait6731;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15585_i\));
                      state_var7021 <= pause_getI6729;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15555_len_aux3143354_result\ := \$15555_len_aux3143354_arg\(36 to 67);
                  \$15455\ := \$15555_len_aux3143354_result\;
                  \$v6727\ := \$$10702_brk_ptr_take\;
                  if \$v6727\(0) = '1' then
                    state_var7021 <= q_wait6726;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6724;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII6759 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15454\ := \$$10699_symtbl_value\;
              \$15555_len_aux3143354_arg\ := \$15240_loop23133355_arg\(0 to 35) & X"0000000" & X"0" & eclat_unit;
              state_var7021 <= \$15555_len_aux3143354\;
            when pause_getII6763 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15319\ := \$$10699_symtbl_value\;
              \$15240_loop23133355_result\ := eclat_unit;
              \$15217_loop1312_result\ := \$15240_loop23133355_result\;
              state_var7021 <= \$14481_decode_loop310\;
            when pause_getII6772 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15317\ := \$$10699_symtbl_value\;
              \$v6770\ := \$$10696_ram_ptr_take\;
              if \$v6770\(0) = '1' then
                state_var7021 <= q_wait6769;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6766\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15317\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15311_end_rib\ & "0000" & \$15293\ & "0001" & \$v6766\;
                state_var7021 <= pause_setI6767;
              end if;
            when pause_getII6780 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15315_i\ := \$$10702_brk_value\;
              \$v6778\ := \$$10699_symtbl_ptr_take\;
              if \$v6778\(0) = '1' then
                state_var7021 <= q_wait6777;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15315_i\;
                state_var7021 <= pause_setI6775;
              end if;
            when pause_getII6784 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15315_i\ := \$$10702_brk_value\;
              \$v6778\ := \$$10699_symtbl_ptr_take\;
              if \$v6778\(0) = '1' then
                state_var7021 <= q_wait6777;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15315_i\;
                state_var7021 <= pause_setI6775;
              end if;
            when pause_getII6792 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15324\ := \$$10702_brk_value\;
              \$v6790\ := \$$10702_brk_ptr_take\;
              if \$v6790\(0) = '1' then
                state_var7021 <= q_wait6789;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15324\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6787;
              end if;
            when pause_getII6797 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15314\ := \$$10695_limit_value\;
              \$v6795\ := eclat_eq(\$15313\ & eclat_sub(\$15314\ & X"0000000" & X"1"));
              if \$v6795\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15332_forever3163343\;
              else
                \$v6794\ := \$$10702_brk_ptr_take\;
                if \$v6794\(0) = '1' then
                  state_var7021 <= q_wait6793;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6791;
                end if;
              end if;
            when pause_getII6801 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15313\ := \$$10702_brk_value\;
              \$v6799\ := \$$10695_limit_ptr_take\;
              if \$v6799\(0) = '1' then
                state_var7021 <= q_wait6798;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6796;
              end if;
            when pause_getII6805 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15342\ := \$$10699_symtbl_value\;
              \$15311_end_rib\ := "0000" & \$15342\;
              \$v6803\ := \$$10702_brk_ptr_take\;
              if \$v6803\(0) = '1' then
                state_var7021 <= q_wait6802;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6800;
              end if;
            when pause_getII6815 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15309\ := \$$10699_symtbl_value\;
              \$v6813\ := \$$10696_ram_ptr_take\;
              if \$v6813\(0) = '1' then
                state_var7021 <= q_wait6812;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6808\ := X"0000000" & X"2";
                \$v6809\ := X"0000000" & X"2";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15309\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v6808\ & \$15303_str_rib\ & "0001" & \$v6809\;
                state_var7021 <= pause_setI6810;
              end if;
            when pause_getII6823 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15307_i\ := \$$10702_brk_value\;
              \$v6821\ := \$$10699_symtbl_ptr_take\;
              if \$v6821\(0) = '1' then
                state_var7021 <= q_wait6820;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15307_i\;
                state_var7021 <= pause_setI6818;
              end if;
            when pause_getII6827 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15307_i\ := \$$10702_brk_value\;
              \$v6821\ := \$$10699_symtbl_ptr_take\;
              if \$v6821\(0) = '1' then
                state_var7021 <= q_wait6820;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15307_i\;
                state_var7021 <= pause_setI6818;
              end if;
            when pause_getII6835 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15347\ := \$$10702_brk_value\;
              \$v6833\ := \$$10702_brk_ptr_take\;
              if \$v6833\(0) = '1' then
                state_var7021 <= q_wait6832;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15347\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6830;
              end if;
            when pause_getII6840 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15306\ := \$$10695_limit_value\;
              \$v6838\ := eclat_eq(\$15305\ & eclat_sub(\$15306\ & X"0000000" & X"1"));
              if \$v6838\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15355_forever3163344\;
              else
                \$v6837\ := \$$10702_brk_ptr_take\;
                if \$v6837\(0) = '1' then
                  state_var7021 <= q_wait6836;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6834;
                end if;
              end if;
            when pause_getII6844 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15305\ := \$$10702_brk_value\;
              \$v6842\ := \$$10695_limit_ptr_take\;
              if \$v6842\(0) = '1' then
                state_var7021 <= q_wait6841;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6839;
              end if;
            when pause_getII6848 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15365\ := \$$10699_symtbl_value\;
              \$15303_str_rib\ := "0000" & \$15365\;
              \$v6846\ := \$$10702_brk_ptr_take\;
              if \$v6846\(0) = '1' then
                state_var7021 <= q_wait6845;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6843;
              end if;
            when pause_getII6857 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15301\ := \$$10699_symtbl_value\;
              \$v6855\ := \$$10696_ram_ptr_take\;
              if \$v6855\(0) = '1' then
                state_var7021 <= q_wait6854;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6851\ := X"0000000" & X"3";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15301\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15240_loop23133355_arg\(0 to 35) & "0001" & \$15294\ & "0001" & \$v6851\;
                state_var7021 <= pause_setI6852;
              end if;
            when pause_getII6865 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15299_i\ := \$$10702_brk_value\;
              \$v6863\ := \$$10699_symtbl_ptr_take\;
              if \$v6863\(0) = '1' then
                state_var7021 <= q_wait6862;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15299_i\;
                state_var7021 <= pause_setI6860;
              end if;
            when pause_getII6869 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15299_i\ := \$$10702_brk_value\;
              \$v6863\ := \$$10699_symtbl_ptr_take\;
              if \$v6863\(0) = '1' then
                state_var7021 <= q_wait6862;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15299_i\;
                state_var7021 <= pause_setI6860;
              end if;
            when pause_getII6877 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15370\ := \$$10702_brk_value\;
              \$v6875\ := \$$10702_brk_ptr_take\;
              if \$v6875\(0) = '1' then
                state_var7021 <= q_wait6874;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15370\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6872;
              end if;
            when pause_getII6882 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15298\ := \$$10695_limit_value\;
              \$v6880\ := eclat_eq(\$15296\ & eclat_sub(\$15298\ & X"0000000" & X"1"));
              if \$v6880\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15378_forever3163345\;
              else
                \$v6879\ := \$$10702_brk_ptr_take\;
                if \$v6879\(0) = '1' then
                  state_var7021 <= q_wait6878;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6876;
                end if;
              end if;
            when pause_getII6886 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15296\ := \$$10702_brk_value\;
              \$v6884\ := \$$10695_limit_ptr_take\;
              if \$v6884\(0) = '1' then
                state_var7021 <= q_wait6883;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6881;
              end if;
            when pause_getII6891 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15401\ := \$$10696_ram_value\;
              \$15391_len_aux3143348_arg\ := \$15401\(36 to 71) & eclat_add(\$15391_len_aux3143348_arg\(36 to 67) & X"0000000" & X"1") & eclat_unit;
              state_var7021 <= \$15391_len_aux3143348\;
            when pause_getII6910 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$15422\ := \$$10696_ram_value\;
              \$v6906\ := \$15422\(72 to 107);
              \$v6907\ := \$v6906\(0 to 3);
              \$v6897\ := \$v6906\(4 to 35);
              case \$v6907\ is
              when "0001" =>
                \$15427_i\ := \$v6897\(0 to 31);
                \$v6901\ := X"0000000" & X"0";
                \$v6899\ := "0001" & \$v6901\;
                \$v6900\ := \$v6899\(0 to 3);
                \$v6898\ := \$v6899\(4 to 35);
                case \$v6900\ is
                when "0000" =>
                  \$15400\ := eclat_false;
                when "0001" =>
                  \$15430_j\ := \$v6898\(0 to 31);
                  \$15400\ := eclat_eq(\$15427_i\ & \$15430_j\);
                when others =>
                  
                end case;
                \$v6896\ := \$15400\;
                if \$v6896\(0) = '1' then
                  \$v6894\ := \$15391_len_aux3143348_arg\(0 to 35);
                  \$v6895\ := \$v6894\(0 to 3);
                  \$v6889\ := \$v6894\(4 to 35);
                  case \$v6895\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15413_forever3163346\;
                  when "0000" =>
                    \$15421_i\ := \$v6889\(0 to 31);
                    \$v6893\ := \$$10696_ram_ptr_take\;
                    if \$v6893\(0) = '1' then
                      state_var7021 <= q_wait6892;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15421_i\));
                      state_var7021 <= pause_getI6890;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15391_len_aux3143348_result\ := \$15391_len_aux3143348_arg\(36 to 67);
                  \$15294\ := \$15391_len_aux3143348_result\;
                  \$v6888\ := \$$10702_brk_ptr_take\;
                  if \$v6888\(0) = '1' then
                    state_var7021 <= q_wait6887;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6885;
                  end if;
                end if;
              when "0000" =>
                \$15431_i\ := \$v6897\(0 to 31);
                \$v6905\ := X"0000000" & X"0";
                \$v6903\ := "0001" & \$v6905\;
                \$v6904\ := \$v6903\(0 to 3);
                \$v6902\ := \$v6903\(4 to 35);
                case \$v6904\ is
                when "0001" =>
                  \$15400\ := eclat_false;
                when "0000" =>
                  \$15434_j\ := \$v6902\(0 to 31);
                  \$15400\ := eclat_eq(\$15431_i\ & \$15434_j\);
                when others =>
                  
                end case;
                \$v6896\ := \$15400\;
                if \$v6896\(0) = '1' then
                  \$v6894\ := \$15391_len_aux3143348_arg\(0 to 35);
                  \$v6895\ := \$v6894\(0 to 3);
                  \$v6889\ := \$v6894\(4 to 35);
                  case \$v6895\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$15413_forever3163346\;
                  when "0000" =>
                    \$15421_i\ := \$v6889\(0 to 31);
                    \$v6893\ := \$$10696_ram_ptr_take\;
                    if \$v6893\(0) = '1' then
                      state_var7021 <= q_wait6892;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$15421_i\));
                      state_var7021 <= pause_getI6890;
                    end if;
                  when others =>
                    
                  end case;
                else
                  \$15391_len_aux3143348_result\ := \$15391_len_aux3143348_arg\(36 to 67);
                  \$15294\ := \$15391_len_aux3143348_result\;
                  \$v6888\ := \$$10702_brk_ptr_take\;
                  if \$v6888\(0) = '1' then
                    state_var7021 <= q_wait6887;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6885;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII6920 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$15293\ := \$$10699_symtbl_value\;
              \$15391_len_aux3143348_arg\ := \$15240_loop23133355_arg\(0 to 35) & X"0000000" & X"0" & eclat_unit;
              state_var7021 <= \$15391_len_aux3143348\;
            when pause_getII6924 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$15268\ := \$$10698_heap_value\;
              \$15267\ := "0000" & \$15268\;
              \$15240_loop23133355_arg\ := \$15267\ & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var7021 <= \$15240_loop23133355\;
            when pause_getII6934 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$15265\ := \$$10698_heap_value\;
              \$v6932\ := \$$10696_ram_ptr_take\;
              if \$v6932\(0) = '1' then
                state_var7021 <= q_wait6931;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6927\ := eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$15255\,32);
                \$v6928\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15265\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v6927\ & \$15240_loop23133355_arg\(0 to 35) & "0001" & \$v6928\;
                state_var7021 <= pause_setI6929;
              end if;
            when pause_getII6942 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15263_i\ := \$$10702_brk_value\;
              \$v6940\ := \$$10698_heap_ptr_take\;
              if \$v6940\(0) = '1' then
                state_var7021 <= q_wait6939;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$15263_i\;
                state_var7021 <= pause_setI6937;
              end if;
            when pause_getII6946 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15263_i\ := \$$10702_brk_value\;
              \$v6940\ := \$$10698_heap_ptr_take\;
              if \$v6940\(0) = '1' then
                state_var7021 <= q_wait6939;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$15263_i\;
                state_var7021 <= pause_setI6937;
              end if;
            when pause_getII6954 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15274\ := \$$10702_brk_value\;
              \$v6952\ := \$$10702_brk_ptr_take\;
              if \$v6952\(0) = '1' then
                state_var7021 <= q_wait6951;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15274\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6949;
              end if;
            when pause_getII6959 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15262\ := \$$10695_limit_value\;
              \$v6957\ := eclat_eq(\$15261\ & eclat_sub(\$15262\ & X"0000000" & X"1"));
              if \$v6957\(0) = '1' then
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not implemented"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$15282_forever3163342\;
              else
                \$v6956\ := \$$10702_brk_ptr_take\;
                if \$v6956\(0) = '1' then
                  state_var7021 <= q_wait6955;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI6953;
                end if;
              end if;
            when pause_getII6963 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$15261\ := \$$10702_brk_value\;
              \$v6961\ := \$$10695_limit_ptr_take\;
              if \$v6961\(0) = '1' then
                state_var7021 <= q_wait6960;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6958;
              end if;
            when pause_getII6973 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$15256\ := \$$10701_pos_value\;
              \$v6971\ := \$$10701_pos_ptr_take\;
              if \$v6971\(0) = '1' then
                state_var7021 <= q_wait6970;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$15256\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6968;
              end if;
            when pause_getII6977 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$15255\ := \$$10701_pos_value\;
              \$v6975\ := \$$10701_pos_ptr_take\;
              if \$v6975\(0) = '1' then
                state_var7021 <= q_wait6974;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6972;
              end if;
            when pause_getII6988 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$15797\ := \$$10701_pos_value\;
              \$v6986\ := \$$10701_pos_ptr_take\;
              if \$v6986\(0) = '1' then
                state_var7021 <= q_wait6985;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$15797\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6983;
              end if;
            when pause_getII6992 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$15796\ := \$$10701_pos_value\;
              \$v6990\ := \$$10701_pos_ptr_take\;
              if \$v6990\(0) = '1' then
                state_var7021 <= q_wait6989;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6987;
              end if;
            when pause_setI3370 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII3371;
            when pause_setI3384 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3385;
            when pause_setI3392 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3393;
            when pause_setI3413 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3414;
            when pause_setI3438 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3439;
            when pause_setI3466 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3467;
            when pause_setI3524 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3525;
            when pause_setI3532 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII3533;
            when pause_setI3544 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII3545;
            when pause_setI3561 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3562;
            when pause_setI3593 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3594;
            when pause_setI3601 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII3602;
            when pause_setI3613 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII3614;
            when pause_setI3630 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII3631;
            when pause_setI3648 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII3649;
            when pause_setI3663 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3664;
            when pause_setI3721 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3722;
            when pause_setI3729 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3730;
            when pause_setI3745 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII3746;
            when pause_setI3766 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3767;
            when pause_setI3774 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII3775;
            when pause_setI3786 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII3787;
            when pause_setI3803 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3804;
            when pause_setI3818 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3819;
            when pause_setI3833 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3834;
            when pause_setI3849 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3850;
            when pause_setI3857 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3858;
            when pause_setI3873 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII3874;
            when pause_setI3890 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3891;
            when pause_setI3905 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3906;
            when pause_setI3921 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3922;
            when pause_setI3929 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3930;
            when pause_setI3945 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII3946;
            when pause_setI3962 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3963;
            when pause_setI3977 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII3978;
            when pause_setI3993 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII3994;
            when pause_setI4001 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4002;
            when pause_setI4017 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4018;
            when pause_setI4039 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4040;
            when pause_setI4047 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII4048;
            when pause_setI4059 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4060;
            when pause_setI4087 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4088;
            when pause_setI4105 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4106;
            when pause_setI4113 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4114;
            when pause_setI4129 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4130;
            when pause_setI4149 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4150;
            when pause_setI4165 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4166;
            when pause_setI4173 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4174;
            when pause_setI4189 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4190;
            when pause_setI4213 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4214;
            when pause_setI4229 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4230;
            when pause_setI4237 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4238;
            when pause_setI4253 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4254;
            when pause_setI4277 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4278;
            when pause_setI4293 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4294;
            when pause_setI4301 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4302;
            when pause_setI4317 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4318;
            when pause_setI4341 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4342;
            when pause_setI4357 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4358;
            when pause_setI4365 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4366;
            when pause_setI4381 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4382;
            when pause_setI4399 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4400;
            when pause_setI4419 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4420;
            when pause_setI4434 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4435;
            when pause_setI4450 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4451;
            when pause_setI4458 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4459;
            when pause_setI4474 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4475;
            when pause_setI4492 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4493;
            when pause_setI4512 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4513;
            when pause_setI4527 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4528;
            when pause_setI4543 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4544;
            when pause_setI4551 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4552;
            when pause_setI4567 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4568;
            when pause_setI4585 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4586;
            when pause_setI4605 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4606;
            when pause_setI4620 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4621;
            when pause_setI4638 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4639;
            when pause_setI4646 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4647;
            when pause_setI4662 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4663;
            when pause_setI4731 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4732;
            when pause_setI4746 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4747;
            when pause_setI4762 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4763;
            when pause_setI4770 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4771;
            when pause_setI4786 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4787;
            when pause_setI4811 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4812;
            when pause_setI4826 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4827;
            when pause_setI4842 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4843;
            when pause_setI4850 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4851;
            when pause_setI4866 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4867;
            when pause_setI4890 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4891;
            when pause_setI4905 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4906;
            when pause_setI4921 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII4922;
            when pause_setI4929 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4930;
            when pause_setI4945 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII4946;
            when pause_setI4969 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4970;
            when pause_setI4984 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII4985;
            when pause_setI5000 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5001;
            when pause_setI5008 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5009;
            when pause_setI5024 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5025;
            when pause_setI5048 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5049;
            when pause_setI5063 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5064;
            when pause_setI5079 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5080;
            when pause_setI5087 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5088;
            when pause_setI5103 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5104;
            when pause_setI5127 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5128;
            when pause_setI5142 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5143;
            when pause_setI5158 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5159;
            when pause_setI5166 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5167;
            when pause_setI5182 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5183;
            when pause_setI5200 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5201;
            when pause_setI5208 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5209;
            when pause_setI5224 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5225;
            when pause_setI5244 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5245;
            when pause_setI5318 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII5319;
            when pause_setI5338 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5339;
            when pause_setI5371 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5372;
            when pause_setI5393 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5394;
            when pause_setI5408 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII5409;
            when pause_setI5427 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5428;
            when pause_setI5435 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5436;
            when pause_setI5451 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5452;
            when pause_setI5497 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII5498;
            when pause_setI5516 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5517;
            when pause_setI5524 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5525;
            when pause_setI5540 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5541;
            when pause_setI5557 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII5558;
            when pause_setI5575 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII5576;
            when pause_setI5594 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5595;
            when pause_setI5623 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII5624;
            when pause_setI5629 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5630;
            when pause_setI5636 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5637;
            when pause_setI5648 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5649;
            when pause_setI5673 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5674;
            when pause_setI5690 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII5691;
            when pause_setI5710 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5711;
            when pause_setI5741 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII5742;
            when pause_setI5761 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5762;
            when pause_setI5792 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII5793;
            when pause_setI5812 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5813;
            when pause_setI5843 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII5844;
            when pause_setI5862 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5863;
            when pause_setI5899 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5900;
            when pause_setI5907 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII5908;
            when pause_setI5919 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII5920;
            when pause_setI5940 =>
              \$$10700_pc_write_request\ <= '0';
              state_var7021 <= pause_setII5941;
            when pause_setI5966 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5967;
            when pause_setI5991 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII5992;
            when pause_setI5999 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII6000;
            when pause_setI6011 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6012;
            when pause_setI6039 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII6040;
            when pause_setI6055 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6056;
            when pause_setI6080 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6081;
            when pause_setI6088 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII6089;
            when pause_setI6100 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6101;
            when pause_setI6142 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6143;
            when pause_setI6150 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII6151;
            when pause_setI6162 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6163;
            when pause_setI6184 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6185;
            when pause_setI6192 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII6193;
            when pause_setI6204 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6205;
            when pause_setI6221 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII6222;
            when pause_setI6237 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6238;
            when pause_setI6262 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6263;
            when pause_setI6270 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII6271;
            when pause_setI6282 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6283;
            when pause_setI6333 =>
              \$$10701_pos_write_request\ <= '0';
              state_var7021 <= pause_setII6334;
            when pause_setI6365 =>
              \$$10701_pos_write_request\ <= '0';
              state_var7021 <= pause_setII6366;
            when pause_setI6381 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6382;
            when pause_setI6389 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII6390;
            when pause_setI6405 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6406;
            when pause_setI6425 =>
              \$$10701_pos_write_request\ <= '0';
              state_var7021 <= pause_setII6426;
            when pause_setI6442 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6443;
            when pause_setI6450 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6451;
            when pause_setI6462 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6463;
            when pause_setI6485 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6486;
            when pause_setI6493 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6494;
            when pause_setI6505 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6506;
            when pause_setI6528 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6529;
            when pause_setI6536 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6537;
            when pause_setI6548 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6549;
            when pause_setI6606 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6607;
            when pause_setI6614 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6615;
            when pause_setI6626 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6627;
            when pause_setI6649 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6650;
            when pause_setI6657 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6658;
            when pause_setI6669 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6670;
            when pause_setI6691 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6692;
            when pause_setI6699 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6700;
            when pause_setI6711 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6712;
            when pause_setI6767 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6768;
            when pause_setI6775 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6776;
            when pause_setI6787 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6788;
            when pause_setI6810 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6811;
            when pause_setI6818 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6819;
            when pause_setI6830 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6831;
            when pause_setI6852 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6853;
            when pause_setI6860 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII6861;
            when pause_setI6872 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6873;
            when pause_setI6929 =>
              \$$10696_ram_write_request\ <= '0';
              state_var7021 <= pause_setII6930;
            when pause_setI6937 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII6938;
            when pause_setI6949 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII6950;
            when pause_setI6968 =>
              \$$10701_pos_write_request\ <= '0';
              state_var7021 <= pause_setII6969;
            when pause_setI6983 =>
              \$$10701_pos_write_request\ <= '0';
              state_var7021 <= pause_setII6984;
            when pause_setI6995 =>
              \$$10695_limit_write_request\ <= '0';
              state_var7021 <= pause_setII6996;
            when pause_setI6999 =>
              \$$10702_brk_write_request\ <= '0';
              state_var7021 <= pause_setII7000;
            when pause_setI7003 =>
              \$$10701_pos_write_request\ <= '0';
              state_var7021 <= pause_setII7004;
            when pause_setI7007 =>
              \$$10699_symtbl_write_request\ <= '0';
              state_var7021 <= pause_setII7008;
            when pause_setI7011 =>
              \$$10698_heap_write_request\ <= '0';
              state_var7021 <= pause_setII7012;
            when pause_setI7015 =>
              \$$10697_stack_write_request\ <= '0';
              state_var7021 <= pause_setII7016;
            when pause_setII3371 =>
              \$$10700_pc_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII3385 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v3382\ := \$10819\(0 to 35);
              \$v3383\ := \$v3382\(0 to 3);
              \$v3377\ := \$v3382\(4 to 35);
              case \$v3383\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10872_forever3163137\;
              when "0000" =>
                \$10880_i\ := \$v3377\(0 to 31);
                \$v3381\ := \$$10696_ram_ptr_take\;
                if \$v3381\(0) = '1' then
                  state_var7021 <= q_wait3380;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$10880_i\));
                  state_var7021 <= pause_getI3378;
                end if;
              when others =>
                
              end case;
            when pause_setII3393 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3389\ := \$10839_s\;
              \$v3390\ := \$v3389\(0 to 3);
              \$v3388\ := \$v3389\(4 to 35);
              case \$v3390\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10885_forever3163138\;
              when "0000" =>
                \$10893_i\ := \$v3388\(0 to 31);
                \$10842\ := \$10893_i\;
                \$v3387\ := \$$10697_stack_ptr_take\;
                if \$v3387\(0) = '1' then
                  state_var7021 <= q_wait3386;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$10842\;
                  state_var7021 <= pause_setI3384;
                end if;
              when others =>
                
              end case;
            when pause_setII3414 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3410\ := \$10828_c2_rib\;
              \$v3411\ := \$v3410\(0 to 3);
              \$v3391\ := \$v3410\(4 to 35);
              case \$v3411\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field2_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11090_forever3163150\;
              when "0000" =>
                \$11098_i\ := \$v3391\(0 to 31);
                \$v3408\ := \$10828_c2_rib\;
                \$v3409\ := \$v3408\(0 to 3);
                \$v3403\ := \$v3408\(4 to 35);
                case \$v3409\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$11126_forever3163152\;
                when "0000" =>
                  \$11134_i\ := \$v3403\(0 to 31);
                  \$v3407\ := \$$10696_ram_ptr_take\;
                  if \$v3407\(0) = '1' then
                    state_var7021 <= q_wait3406;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$11134_i\));
                    state_var7021 <= pause_getI3404;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_setII3439 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3389\ := \$10839_s\;
              \$v3390\ := \$v3389\(0 to 3);
              \$v3388\ := \$v3389\(4 to 35);
              case \$v3390\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't int_of_triplet"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10885_forever3163138\;
              when "0000" =>
                \$10893_i\ := \$v3388\(0 to 31);
                \$10842\ := \$10893_i\;
                \$v3387\ := \$$10697_stack_ptr_take\;
                if \$v3387\(0) = '1' then
                  state_var7021 <= q_wait3386;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr_write\ <= 0;
                  \$$10697_stack_write_request\ <= '1';
                  \$$10697_stack_write\ <= \$10842\;
                  state_var7021 <= pause_setI3384;
                end if;
              when others =>
                
              end case;
            when pause_setII3467 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3463\ := \$10897_k\;
              \$v3464\ := \$v3463\(0 to 3);
              \$v3458\ := \$v3463\(4 to 35);
              case \$v3464\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$10958_forever3163142\;
              when "0000" =>
                \$10966_i\ := \$v3458\(0 to 31);
                \$v3462\ := \$$10696_ram_ptr_take\;
                if \$v3462\(0) = '1' then
                  state_var7021 <= q_wait3461;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$10966_i\));
                  state_var7021 <= pause_getI3459;
                end if;
              when others =>
                
              end case;
            when pause_setII3525 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3522\ := \$$10698_heap_ptr_take\;
              if \$v3522\(0) = '1' then
                state_var7021 <= q_wait3521;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3519;
              end if;
            when pause_setII3533 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v3531\ := \$$10698_heap_ptr_take\;
              if \$v3531\(0) = '1' then
                state_var7021 <= q_wait3530;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3528;
              end if;
            when pause_setII3545 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v3543\ := \$$10702_brk_ptr_take\;
              if \$v3543\(0) = '1' then
                state_var7021 <= q_wait3542;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3540;
              end if;
            when pause_setII3562 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11219\ := \$11214\(0 to 35);
              \$v3560\ := \$$10702_brk_ptr_take\;
              if \$v3560\(0) = '1' then
                state_var7021 <= q_wait3559;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3557;
              end if;
            when pause_setII3594 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3590\ := \$$10698_heap_ptr_take\;
              if \$v3590\(0) = '1' then
                state_var7021 <= q_wait3589;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3587;
              end if;
            when pause_setII3602 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v3600\ := \$$10698_heap_ptr_take\;
              if \$v3600\(0) = '1' then
                state_var7021 <= q_wait3599;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3597;
              end if;
            when pause_setII3614 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v3612\ := \$$10702_brk_ptr_take\;
              if \$v3612\(0) = '1' then
                state_var7021 <= q_wait3611;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3609;
              end if;
            when pause_setII3631 =>
              \$$10700_pc_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII3649 =>
              \$$10700_pc_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII3664 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3660\ := \$11328_cont\;
              \$v3661\ := \$v3660\(0 to 3);
              \$v3655\ := \$v3660\(4 to 35);
              case \$v3661\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11356_forever3163163\;
              when "0000" =>
                \$11364_i\ := \$v3655\(0 to 31);
                \$v3659\ := \$$10696_ram_ptr_take\;
                if \$v3659\(0) = '1' then
                  state_var7021 <= q_wait3658;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11364_i\));
                  state_var7021 <= pause_getI3656;
                end if;
              when others =>
                
              end case;
            when pause_setII3722 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII3730 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v3728\ := \$$10697_stack_ptr_take\;
              if \$v3728\(0) = '1' then
                state_var7021 <= q_wait3727;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3725;
              end if;
            when pause_setII3746 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v3744\ := \$$10702_brk_ptr_take\;
              if \$v3744\(0) = '1' then
                state_var7021 <= q_wait3743;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3741;
              end if;
            when pause_setII3767 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3765\ := \$$10698_heap_ptr_take\;
              if \$v3765\(0) = '1' then
                state_var7021 <= q_wait3764;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3762;
              end if;
            when pause_setII3775 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v3773\ := \$$10698_heap_ptr_take\;
              if \$v3773\(0) = '1' then
                state_var7021 <= q_wait3772;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3770;
              end if;
            when pause_setII3787 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v3785\ := \$$10702_brk_ptr_take\;
              if \$v3785\(0) = '1' then
                state_var7021 <= q_wait3784;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3782;
              end if;
            when pause_setII3804 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11556_z\ := \$11551\(0 to 35);
              \$v3802\ := \$$10702_brk_ptr_take\;
              if \$v3802\(0) = '1' then
                state_var7021 <= q_wait3801;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3799;
              end if;
            when pause_setII3819 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11548_y\ := \$11543\(0 to 35);
              \$v3817\ := \$$10697_stack_ptr_take\;
              if \$v3817\(0) = '1' then
                state_var7021 <= q_wait3816;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3814;
              end if;
            when pause_setII3834 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11540_x\ := \$11535\(0 to 35);
              \$v3832\ := \$$10697_stack_ptr_take\;
              if \$v3832\(0) = '1' then
                state_var7021 <= q_wait3831;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3829;
              end if;
            when pause_setII3850 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII3858 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v3856\ := \$$10697_stack_ptr_take\;
              if \$v3856\(0) = '1' then
                state_var7021 <= q_wait3855;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3853;
              end if;
            when pause_setII3874 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v3872\ := \$$10702_brk_ptr_take\;
              if \$v3872\(0) = '1' then
                state_var7021 <= q_wait3871;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3869;
              end if;
            when pause_setII3891 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11663\ := \$11658\(0 to 35);
              \$v3889\ := \$$10702_brk_ptr_take\;
              if \$v3889\(0) = '1' then
                state_var7021 <= q_wait3888;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3886;
              end if;
            when pause_setII3906 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII3922 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII3930 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v3928\ := \$$10697_stack_ptr_take\;
              if \$v3928\(0) = '1' then
                state_var7021 <= q_wait3927;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3925;
              end if;
            when pause_setII3946 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v3944\ := \$$10702_brk_ptr_take\;
              if \$v3944\(0) = '1' then
                state_var7021 <= q_wait3943;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3941;
              end if;
            when pause_setII3963 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v3961\ := \$$10702_brk_ptr_take\;
              if \$v3961\(0) = '1' then
                state_var7021 <= q_wait3960;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3958;
              end if;
            when pause_setII3978 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11736_x\ := \$11731\(0 to 35);
              \$v3976\ := \$$10697_stack_ptr_take\;
              if \$v3976\(0) = '1' then
                state_var7021 <= q_wait3975;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3973;
              end if;
            when pause_setII3994 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4002 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4000\ := \$$10697_stack_ptr_take\;
              if \$v4000\(0) = '1' then
                state_var7021 <= q_wait3999;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3997;
              end if;
            when pause_setII4018 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4016\ := \$$10702_brk_ptr_take\;
              if \$v4016\(0) = '1' then
                state_var7021 <= q_wait4015;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4013;
              end if;
            when pause_setII4040 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v4037\ := \$$10698_heap_ptr_take\;
              if \$v4037\(0) = '1' then
                state_var7021 <= q_wait4036;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI4034;
              end if;
            when pause_setII4048 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v4046\ := \$$10698_heap_ptr_take\;
              if \$v4046\(0) = '1' then
                state_var7021 <= q_wait4045;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI4043;
              end if;
            when pause_setII4060 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4058\ := \$$10702_brk_ptr_take\;
              if \$v4058\(0) = '1' then
                state_var7021 <= q_wait4057;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4055;
              end if;
            when pause_setII4088 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11809\ := \$11804\(0 to 35);
              \$v4085\ := \$11809\;
              \$v4086\ := \$v4085\(0 to 3);
              \$v4080\ := \$v4085\(4 to 35);
              case \$v4086\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$11881_forever3163187\;
              when "0000" =>
                \$11889_i\ := \$v4080\(0 to 31);
                \$v4084\ := \$$10696_ram_ptr_take\;
                if \$v4084\(0) = '1' then
                  state_var7021 <= q_wait4083;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$11889_i\));
                  state_var7021 <= pause_getI4081;
                end if;
              when others =>
                
              end case;
            when pause_setII4106 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4114 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4112\ := \$$10697_stack_ptr_take\;
              if \$v4112\(0) = '1' then
                state_var7021 <= q_wait4111;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4109;
              end if;
            when pause_setII4130 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4128\ := \$$10702_brk_ptr_take\;
              if \$v4128\(0) = '1' then
                state_var7021 <= q_wait4127;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4125;
              end if;
            when pause_setII4150 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11911\ := \$11906\(0 to 35);
              \$v4147\ := \$11911\;
              \$v4148\ := \$v4147\(0 to 3);
              \$v4146\ := \$v4147\(4 to 35);
              case \$v4148\ is
              when "0001" =>
                \$11912\ := eclat_false;
              when "0000" =>
                \$11944_i\ := \$v4146\(0 to 31);
                \$11912\ := eclat_if(eclat_ge(\$11944_i\ & X"0000000" & X"0") & eclat_lt(\$11944_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v4145\ := \$$10702_brk_ptr_take\;
              if \$v4145\(0) = '1' then
                state_var7021 <= q_wait4144;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4142;
              end if;
            when pause_setII4166 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4174 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4172\ := \$$10697_stack_ptr_take\;
              if \$v4172\(0) = '1' then
                state_var7021 <= q_wait4171;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4169;
              end if;
            when pause_setII4190 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4188\ := \$$10702_brk_ptr_take\;
              if \$v4188\(0) = '1' then
                state_var7021 <= q_wait4187;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4185;
              end if;
            when pause_setII4214 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$11967\ := \$11962\(0 to 35);
              \$v4211\ := \$11967\;
              \$v4212\ := \$v4211\(0 to 3);
              \$v4206\ := \$v4211\(4 to 35);
              case \$v4212\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12006_forever3163192\;
              when "0000" =>
                \$12014_i\ := \$v4206\(0 to 31);
                \$v4210\ := \$$10696_ram_ptr_take\;
                if \$v4210\(0) = '1' then
                  state_var7021 <= q_wait4209;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$12014_i\));
                  state_var7021 <= pause_getI4207;
                end if;
              when others =>
                
              end case;
            when pause_setII4230 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4238 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4236\ := \$$10697_stack_ptr_take\;
              if \$v4236\(0) = '1' then
                state_var7021 <= q_wait4235;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4233;
              end if;
            when pause_setII4254 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4252\ := \$$10702_brk_ptr_take\;
              if \$v4252\(0) = '1' then
                state_var7021 <= q_wait4251;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4249;
              end if;
            when pause_setII4278 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12036\ := \$12031\(0 to 35);
              \$v4275\ := \$12036\;
              \$v4276\ := \$v4275\(0 to 3);
              \$v4270\ := \$v4275\(4 to 35);
              case \$v4276\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12075_forever3163195\;
              when "0000" =>
                \$12083_i\ := \$v4270\(0 to 31);
                \$v4274\ := \$$10696_ram_ptr_take\;
                if \$v4274\(0) = '1' then
                  state_var7021 <= q_wait4273;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$12083_i\));
                  state_var7021 <= pause_getI4271;
                end if;
              when others =>
                
              end case;
            when pause_setII4294 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4302 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4300\ := \$$10697_stack_ptr_take\;
              if \$v4300\(0) = '1' then
                state_var7021 <= q_wait4299;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4297;
              end if;
            when pause_setII4318 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4316\ := \$$10702_brk_ptr_take\;
              if \$v4316\(0) = '1' then
                state_var7021 <= q_wait4315;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4313;
              end if;
            when pause_setII4342 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12105\ := \$12100\(0 to 35);
              \$v4339\ := \$12105\;
              \$v4340\ := \$v4339\(0 to 3);
              \$v4334\ := \$v4339\(4 to 35);
              case \$v4340\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't get_rib"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12144_forever3163198\;
              when "0000" =>
                \$12152_i\ := \$v4334\(0 to 31);
                \$v4338\ := \$$10696_ram_ptr_take\;
                if \$v4338\(0) = '1' then
                  state_var7021 <= q_wait4337;
                else
                  \$$10696_ram_ptr_take\(0) := '1';
                  \$$10696_ram_ptr\ <= to_integer(unsigned(\$12152_i\));
                  state_var7021 <= pause_getI4335;
                end if;
              when others =>
                
              end case;
            when pause_setII4358 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4366 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4364\ := \$$10697_stack_ptr_take\;
              if \$v4364\(0) = '1' then
                state_var7021 <= q_wait4363;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4361;
              end if;
            when pause_setII4382 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4380\ := \$$10702_brk_ptr_take\;
              if \$v4380\(0) = '1' then
                state_var7021 <= q_wait4379;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4377;
              end if;
            when pause_setII4400 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v4397\ := \$$10702_brk_ptr_take\;
              if \$v4397\(0) = '1' then
                state_var7021 <= q_wait4396;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4394;
              end if;
            when pause_setII4420 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12182_y\ := \$12177\(0 to 35);
              \$v4417\ := \$12182_y\;
              \$v4418\ := \$v4417\(0 to 3);
              \$v4398\ := \$v4417\(4 to 35);
              case \$v4418\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field0_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12217_forever3163201\;
              when "0000" =>
                \$12225_i\ := \$v4398\(0 to 31);
                \$v4415\ := \$12182_y\;
                \$v4416\ := \$v4415\(0 to 3);
                \$v4410\ := \$v4415\(4 to 35);
                case \$v4416\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$12253_forever3163203\;
                when "0000" =>
                  \$12261_i\ := \$v4410\(0 to 31);
                  \$v4414\ := \$$10696_ram_ptr_take\;
                  if \$v4414\(0) = '1' then
                    state_var7021 <= q_wait4413;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$12261_i\));
                    state_var7021 <= pause_getI4411;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_setII4435 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12174_x\ := \$12169\(0 to 35);
              \$v4433\ := \$$10697_stack_ptr_take\;
              if \$v4433\(0) = '1' then
                state_var7021 <= q_wait4432;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4430;
              end if;
            when pause_setII4451 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4459 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4457\ := \$$10697_stack_ptr_take\;
              if \$v4457\(0) = '1' then
                state_var7021 <= q_wait4456;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4454;
              end if;
            when pause_setII4475 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4473\ := \$$10702_brk_ptr_take\;
              if \$v4473\(0) = '1' then
                state_var7021 <= q_wait4472;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4470;
              end if;
            when pause_setII4493 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v4490\ := \$$10702_brk_ptr_take\;
              if \$v4490\(0) = '1' then
                state_var7021 <= q_wait4489;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4487;
              end if;
            when pause_setII4513 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12305_y\ := \$12300\(0 to 35);
              \$v4510\ := \$12305_y\;
              \$v4511\ := \$v4510\(0 to 3);
              \$v4491\ := \$v4510\(4 to 35);
              case \$v4511\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field1_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12340_forever3163207\;
              when "0000" =>
                \$12348_i\ := \$v4491\(0 to 31);
                \$v4508\ := \$12305_y\;
                \$v4509\ := \$v4508\(0 to 3);
                \$v4503\ := \$v4508\(4 to 35);
                case \$v4509\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$12376_forever3163209\;
                when "0000" =>
                  \$12384_i\ := \$v4503\(0 to 31);
                  \$v4507\ := \$$10696_ram_ptr_take\;
                  if \$v4507\(0) = '1' then
                    state_var7021 <= q_wait4506;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$12384_i\));
                    state_var7021 <= pause_getI4504;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_setII4528 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12297_x\ := \$12292\(0 to 35);
              \$v4526\ := \$$10697_stack_ptr_take\;
              if \$v4526\(0) = '1' then
                state_var7021 <= q_wait4525;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4523;
              end if;
            when pause_setII4544 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4552 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4550\ := \$$10697_stack_ptr_take\;
              if \$v4550\(0) = '1' then
                state_var7021 <= q_wait4549;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4547;
              end if;
            when pause_setII4568 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4566\ := \$$10702_brk_ptr_take\;
              if \$v4566\(0) = '1' then
                state_var7021 <= q_wait4565;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4563;
              end if;
            when pause_setII4586 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v4583\ := \$$10702_brk_ptr_take\;
              if \$v4583\(0) = '1' then
                state_var7021 <= q_wait4582;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4580;
              end if;
            when pause_setII4606 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12428_y\ := \$12423\(0 to 35);
              \$v4603\ := \$12428_y\;
              \$v4604\ := \$v4603\(0 to 3);
              \$v4584\ := \$v4603\(4 to 35);
              case \$v4604\ is
              when "0001" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't field2_set"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12463_forever3163213\;
              when "0000" =>
                \$12471_i\ := \$v4584\(0 to 31);
                \$v4601\ := \$12428_y\;
                \$v4602\ := \$v4601\(0 to 3);
                \$v4596\ := \$v4601\(4 to 35);
                case \$v4602\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't get_rib"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$12499_forever3163215\;
                when "0000" =>
                  \$12507_i\ := \$v4596\(0 to 31);
                  \$v4600\ := \$$10696_ram_ptr_take\;
                  if \$v4600\(0) = '1' then
                    state_var7021 <= q_wait4599;
                  else
                    \$$10696_ram_ptr_take\(0) := '1';
                    \$$10696_ram_ptr\ <= to_integer(unsigned(\$12507_i\));
                    state_var7021 <= pause_getI4597;
                  end if;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_setII4621 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12420_x\ := \$12415\(0 to 35);
              \$v4619\ := \$$10697_stack_ptr_take\;
              if \$v4619\(0) = '1' then
                state_var7021 <= q_wait4618;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4616;
              end if;
            when pause_setII4639 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4647 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4645\ := \$$10697_stack_ptr_take\;
              if \$v4645\(0) = '1' then
                state_var7021 <= q_wait4644;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4642;
              end if;
            when pause_setII4663 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4661\ := \$$10702_brk_ptr_take\;
              if \$v4661\(0) = '1' then
                state_var7021 <= q_wait4660;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4658;
              end if;
            when pause_setII4732 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12551_y\ := \$12546\(0 to 35);
              \$v4729\ := \$12551_y\;
              \$v4730\ := \$v4729\(0 to 3);
              \$v4679\ := \$v4729\(4 to 35);
              case \$v4730\ is
              when "0001" =>
                \$12583_i\ := \$v4679\(0 to 31);
                \$v4681\ := \$12543_x\;
                \$v4682\ := \$v4681\(0 to 3);
                \$v4680\ := \$v4681\(4 to 35);
                case \$v4682\ is
                when "0001" =>
                  \$12584_j\ := \$v4680\(0 to 31);
                  \$12552\ := eclat_eq(\$12583_i\ & \$12584_j\);
                when others =>
                  \$12552\ := eclat_false;
                end case;
                \$v4678\ := \$$10702_brk_ptr_take\;
                if \$v4678\(0) = '1' then
                  state_var7021 <= q_wait4677;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI4675;
                end if;
              when "0000" =>
                \$v4727\ := \$12543_x\;
                \$v4728\ := \$v4727\(0 to 3);
                \$v4683\ := \$v4727\(4 to 35);
                case \$v4728\ is
                when "0000" =>
                  \$v4725\ := \$12551_y\;
                  \$v4726\ := \$v4725\(0 to 3);
                  \$v4720\ := \$v4725\(4 to 35);
                  case \$v4726\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$12634_forever3163220\;
                  when "0000" =>
                    \$12642_i\ := \$v4720\(0 to 31);
                    \$v4724\ := \$$10696_ram_ptr_take\;
                    if \$v4724\(0) = '1' then
                      state_var7021 <= q_wait4723;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$12642_i\));
                      state_var7021 <= pause_getI4721;
                    end if;
                  when others =>
                    
                  end case;
                when others =>
                  \$12552\ := eclat_false;
                  \$v4678\ := \$$10702_brk_ptr_take\;
                  if \$v4678\(0) = '1' then
                    state_var7021 <= q_wait4677;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI4675;
                  end if;
                end case;
              when others =>
                
              end case;
            when pause_setII4747 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12543_x\ := \$12538\(0 to 35);
              \$v4745\ := \$$10697_stack_ptr_take\;
              if \$v4745\(0) = '1' then
                state_var7021 <= q_wait4744;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4742;
              end if;
            when pause_setII4763 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4771 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4769\ := \$$10697_stack_ptr_take\;
              if \$v4769\(0) = '1' then
                state_var7021 <= q_wait4768;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4766;
              end if;
            when pause_setII4787 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4785\ := \$$10702_brk_ptr_take\;
              if \$v4785\(0) = '1' then
                state_var7021 <= q_wait4784;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4782;
              end if;
            when pause_setII4812 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12686_y\ := \$12681\(0 to 35);
              \$v4809\ := \$12678_x\;
              \$v4810\ := \$v4809\(0 to 3);
              \$v4803\ := \$v4809\(4 to 35);
              case \$v4810\ is
              when "0001" =>
                \$12717_b\ := \$v4803\(0 to 31);
                \$v4807\ := \$12686_y\;
                \$v4808\ := \$v4807\(0 to 3);
                \$v4804\ := \$v4807\(4 to 35);
                case \$v4808\ is
                when "0001" =>
                  \$12718_a\ := \$v4804\(0 to 31);
                  \$v4806\ := X"0000000" & X"1";
                  \$v4805\ := X"0000000" & X"2";
                  \$12687\ := eclat_if(eclat_lt(\$12718_a\ & \$12717_b\) & "0000" & \$v4806\ & "0000" & \$v4805\);
                  \$v4802\ := \$$10702_brk_ptr_take\;
                  if \$v4802\(0) = '1' then
                    state_var7021 <= q_wait4801;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI4799;
                  end if;
                when others =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("not integer"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$12723_forever3163225\;
                end case;
              when others =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not integer"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12734_forever3163224\;
              end case;
            when pause_setII4827 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12678_x\ := \$12673\(0 to 35);
              \$v4825\ := \$$10697_stack_ptr_take\;
              if \$v4825\(0) = '1' then
                state_var7021 <= q_wait4824;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4822;
              end if;
            when pause_setII4843 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4851 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4849\ := \$$10697_stack_ptr_take\;
              if \$v4849\(0) = '1' then
                state_var7021 <= q_wait4848;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4846;
              end if;
            when pause_setII4867 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4865\ := \$$10702_brk_ptr_take\;
              if \$v4865\(0) = '1' then
                state_var7021 <= q_wait4864;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4862;
              end if;
            when pause_setII4891 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12785_y\ := \$12780\(0 to 35);
              \$v4888\ := \$12777_x\;
              \$v4889\ := \$v4888\(0 to 3);
              \$v4883\ := \$v4888\(4 to 35);
              case \$v4889\ is
              when "0000" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not integer"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12820_forever3163229\;
              when "0001" =>
                \$12828_b\ := \$v4883\(0 to 31);
                \$v4886\ := \$12785_y\;
                \$v4887\ := \$v4886\(0 to 3);
                \$v4884\ := \$v4886\(4 to 35);
                case \$v4887\ is
                when "0001" =>
                  \$12829_a\ := \$v4884\(0 to 31);
                  \$v4885\ := eclat_add(\$12829_a\ & \$12828_b\);
                  \$12786\ := "0001" & \$v4885\;
                  \$v4882\ := \$$10702_brk_ptr_take\;
                  if \$v4882\(0) = '1' then
                    state_var7021 <= q_wait4881;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI4879;
                  end if;
                when others =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("not integer"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$12834_forever3163230\;
                end case;
              when others =>
                
              end case;
            when pause_setII4906 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12777_x\ := \$12772\(0 to 35);
              \$v4904\ := \$$10697_stack_ptr_take\;
              if \$v4904\(0) = '1' then
                state_var7021 <= q_wait4903;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4901;
              end if;
            when pause_setII4922 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII4930 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v4928\ := \$$10697_stack_ptr_take\;
              if \$v4928\(0) = '1' then
                state_var7021 <= q_wait4927;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4925;
              end if;
            when pause_setII4946 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v4944\ := \$$10702_brk_ptr_take\;
              if \$v4944\(0) = '1' then
                state_var7021 <= q_wait4943;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4941;
              end if;
            when pause_setII4970 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12885_y\ := \$12880\(0 to 35);
              \$v4967\ := \$12877_x\;
              \$v4968\ := \$v4967\(0 to 3);
              \$v4962\ := \$v4967\(4 to 35);
              case \$v4968\ is
              when "0000" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not integer"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$12920_forever3163234\;
              when "0001" =>
                \$12928_b\ := \$v4962\(0 to 31);
                \$v4965\ := \$12885_y\;
                \$v4966\ := \$v4965\(0 to 3);
                \$v4963\ := \$v4965\(4 to 35);
                case \$v4966\ is
                when "0001" =>
                  \$12929_a\ := \$v4963\(0 to 31);
                  \$v4964\ := eclat_sub(\$12929_a\ & \$12928_b\);
                  \$12886\ := "0001" & \$v4964\;
                  \$v4961\ := \$$10702_brk_ptr_take\;
                  if \$v4961\(0) = '1' then
                    state_var7021 <= q_wait4960;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI4958;
                  end if;
                when others =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("not integer"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$12934_forever3163235\;
                end case;
              when others =>
                
              end case;
            when pause_setII4985 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12877_x\ := \$12872\(0 to 35);
              \$v4983\ := \$$10697_stack_ptr_take\;
              if \$v4983\(0) = '1' then
                state_var7021 <= q_wait4982;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4980;
              end if;
            when pause_setII5001 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII5009 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v5007\ := \$$10697_stack_ptr_take\;
              if \$v5007\(0) = '1' then
                state_var7021 <= q_wait5006;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5004;
              end if;
            when pause_setII5025 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5023\ := \$$10702_brk_ptr_take\;
              if \$v5023\(0) = '1' then
                state_var7021 <= q_wait5022;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5020;
              end if;
            when pause_setII5049 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12985_y\ := \$12980\(0 to 35);
              \$v5046\ := \$12977_x\;
              \$v5047\ := \$v5046\(0 to 3);
              \$v5041\ := \$v5046\(4 to 35);
              case \$v5047\ is
              when "0000" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not integer"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13020_forever3163239\;
              when "0001" =>
                \$13028_b\ := \$v5041\(0 to 31);
                \$v5044\ := \$12985_y\;
                \$v5045\ := \$v5044\(0 to 3);
                \$v5042\ := \$v5044\(4 to 35);
                case \$v5045\ is
                when "0001" =>
                  \$13029_a\ := \$v5042\(0 to 31);
                  \$v5043\ := eclat_mult(\$13029_a\ & \$13028_b\);
                  \$12986\ := "0001" & \$v5043\;
                  \$v5040\ := \$$10702_brk_ptr_take\;
                  if \$v5040\(0) = '1' then
                    state_var7021 <= q_wait5039;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI5037;
                  end if;
                when others =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("not integer"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13034_forever3163240\;
                end case;
              when others =>
                
              end case;
            when pause_setII5064 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$12977_x\ := \$12972\(0 to 35);
              \$v5062\ := \$$10697_stack_ptr_take\;
              if \$v5062\(0) = '1' then
                state_var7021 <= q_wait5061;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5059;
              end if;
            when pause_setII5080 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII5088 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v5086\ := \$$10697_stack_ptr_take\;
              if \$v5086\(0) = '1' then
                state_var7021 <= q_wait5085;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5083;
              end if;
            when pause_setII5104 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5102\ := \$$10702_brk_ptr_take\;
              if \$v5102\(0) = '1' then
                state_var7021 <= q_wait5101;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5099;
              end if;
            when pause_setII5128 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13085_y\ := \$13080\(0 to 35);
              \$v5125\ := \$13077_x\;
              \$v5126\ := \$v5125\(0 to 3);
              \$v5120\ := \$v5125\(4 to 35);
              case \$v5126\ is
              when "0000" =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("not integer"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13120_forever3163244\;
              when "0001" =>
                \$13128_b\ := \$v5120\(0 to 31);
                \$v5123\ := \$13085_y\;
                \$v5124\ := \$v5123\(0 to 3);
                \$v5121\ := \$v5123\(4 to 35);
                case \$v5124\ is
                when "0001" =>
                  \$13129_a\ := \$v5121\(0 to 31);
                  \$v5122\ := eclat_div(\$13129_a\ & \$13128_b\);
                  \$13086\ := "0001" & \$v5122\;
                  \$v5119\ := \$$10702_brk_ptr_take\;
                  if \$v5119\(0) = '1' then
                    state_var7021 <= q_wait5118;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI5116;
                  end if;
                when others =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("not integer"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13134_forever3163245\;
                end case;
              when others =>
                
              end case;
            when pause_setII5143 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13077_x\ := \$13072\(0 to 35);
              \$v5141\ := \$$10697_stack_ptr_take\;
              if \$v5141\(0) = '1' then
                state_var7021 <= q_wait5140;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5138;
              end if;
            when pause_setII5159 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII5167 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v5165\ := \$$10697_stack_ptr_take\;
              if \$v5165\(0) = '1' then
                state_var7021 <= q_wait5164;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5162;
              end if;
            when pause_setII5183 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5181\ := \$$10702_brk_ptr_take\;
              if \$v5181\(0) = '1' then
                state_var7021 <= q_wait5180;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5178;
              end if;
            when pause_setII5201 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v3718\ := \$10814\(72 to 107);
              \$v3719\ := \$v3718\(0 to 3);
              \$v3717\ := \$v3718\(4 to 35);
              case \$v3719\ is
              when "0001" =>
                \$11323\ := eclat_false;
              when "0000" =>
                \$11520_i\ := \$v3717\(0 to 31);
                \$11323\ := eclat_if(eclat_ge(\$11520_i\ & X"0000000" & X"0") & eclat_lt(\$11520_i\ & X"0000" & X"2710") & eclat_false);
              when others =>
                
              end case;
              \$v3716\ := \$11323\;
              if \$v3716\(0) = '1' then
                \$v3647\ := \$$10700_pc_ptr_take\;
                if \$v3647\(0) = '1' then
                  state_var7021 <= q_wait3646;
                else
                  \$$10700_pc_ptr_take\(0) := '1';
                  \$$10700_pc_ptr\ <= 0;
                  state_var7021 <= pause_getI3644;
                end if;
              else
                \$v3715\ := \$$10697_stack_ptr_take\;
                if \$v3715\(0) = '1' then
                  state_var7021 <= q_wait3714;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI3712;
                end if;
              end if;
            when pause_setII5209 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v5207\ := \$$10697_stack_ptr_take\;
              if \$v5207\(0) = '1' then
                state_var7021 <= q_wait5206;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5204;
              end if;
            when pause_setII5225 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5223\ := \$$10702_brk_ptr_take\;
              if \$v5223\(0) = '1' then
                state_var7021 <= q_wait5222;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5220;
              end if;
            when pause_setII5245 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13221\ := \$13216\(0 to 35);
              \$v5242\ := \$13221\;
              \$v5243\ := \$v5242\(0 to 3);
              \$v5241\ := \$v5242\(4 to 35);
              case \$v5243\ is
              when "0001" =>
                \$13252_c\ := \$v5241\(0 to 31);
                eclat_print_char(\$13252_c\);
                
                \$13222\ := "0001" & \$13252_c\;
                \$v5240\ := \$$10702_brk_ptr_take\;
                if \$v5240\(0) = '1' then
                  state_var7021 <= q_wait5239;
                else
                  \$$10702_brk_ptr_take\(0) := '1';
                  \$$10702_brk_ptr\ <= 0;
                  state_var7021 <= pause_getI5237;
                end if;
              when others =>
                eclat_print_string(of_string("Fatal error : "));
                
                eclat_print_string(of_string("can't putchar_prim"));
                
                eclat_print_newline(eclat_unit);
                
                state_var7021 <= \$13257_forever3163251\;
              end case;
            when pause_setII5319 =>
              \$$10700_pc_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII5339 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5335\ := \$$10700_pc_ptr_take\;
              if \$v5335\(0) = '1' then
                state_var7021 <= q_wait5334;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5332;
              end if;
            when pause_setII5372 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5335\ := \$$10700_pc_ptr_take\;
              if \$v5335\(0) = '1' then
                state_var7021 <= q_wait5334;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5332;
              end if;
            when pause_setII5394 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13405\ := \$13400\(0 to 35);
              \$v5391\ := \$10793\(36 to 71);
              \$v5392\ := \$v5391\(0 to 3);
              \$v5336\ := \$v5391\(4 to 35);
              case \$v5392\ is
              when "0001" =>
                \$13443_i\ := \$v5336\(0 to 31);
                \$v5369\ := \$$10697_stack_ptr_take\;
                if \$v5369\(0) = '1' then
                  state_var7021 <= q_wait5368;
                else
                  \$$10697_stack_ptr_take\(0) := '1';
                  \$$10697_stack_ptr\ <= 0;
                  state_var7021 <= pause_getI5366;
                end if;
              when "0000" =>
                \$v5389\ := \$10793\(36 to 71);
                \$v5390\ := \$v5389\(0 to 3);
                \$v5370\ := \$v5389\(4 to 35);
                case \$v5390\ is
                when "0001" =>
                  eclat_print_string(of_string("Fatal error : "));
                  
                  eclat_print_string(of_string("can't field0_set"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var7021 <= \$13537_forever3163267\;
                when "0000" =>
                  \$13545_i\ := \$v5370\(0 to 31);
                  \$v5387\ := \$10793\(36 to 71);
                  \$v5388\ := \$v5387\(0 to 3);
                  \$v5382\ := \$v5387\(4 to 35);
                  case \$v5388\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't get_rib"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$13573_forever3163269\;
                  when "0000" =>
                    \$13581_i\ := \$v5382\(0 to 31);
                    \$v5386\ := \$$10696_ram_ptr_take\;
                    if \$v5386\(0) = '1' then
                      state_var7021 <= q_wait5385;
                    else
                      \$$10696_ram_ptr_take\(0) := '1';
                      \$$10696_ram_ptr\ <= to_integer(unsigned(\$13581_i\));
                      state_var7021 <= pause_getI5383;
                    end if;
                  when others =>
                    
                  end case;
                when others =>
                  
                end case;
              when others =>
                
              end case;
            when pause_setII5409 =>
              \$$10700_pc_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII5428 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5425\ := \$$10700_pc_ptr_take\;
              if \$v5425\(0) = '1' then
                state_var7021 <= q_wait5424;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5422;
              end if;
            when pause_setII5436 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v5434\ := \$$10697_stack_ptr_take\;
              if \$v5434\(0) = '1' then
                state_var7021 <= q_wait5433;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5431;
              end if;
            when pause_setII5452 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5450\ := \$$10702_brk_ptr_take\;
              if \$v5450\(0) = '1' then
                state_var7021 <= q_wait5449;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5447;
              end if;
            when pause_setII5498 =>
              \$$10700_pc_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII5517 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5514\ := \$$10700_pc_ptr_take\;
              if \$v5514\(0) = '1' then
                state_var7021 <= q_wait5513;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5511;
              end if;
            when pause_setII5525 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v5523\ := \$$10697_stack_ptr_take\;
              if \$v5523\(0) = '1' then
                state_var7021 <= q_wait5522;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5520;
              end if;
            when pause_setII5541 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5539\ := \$$10702_brk_ptr_take\;
              if \$v5539\(0) = '1' then
                state_var7021 <= q_wait5538;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5536;
              end if;
            when pause_setII5558 =>
              \$$10700_pc_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII5576 =>
              \$$10700_pc_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII5595 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$13813\ := \$13808\(0 to 35);
              \$v5592\ := \$13813\;
              \$v5593\ := \$v5592\(0 to 3);
              \$v5583\ := \$v5592\(4 to 35);
              case \$v5593\ is
              when "0001" =>
                \$13865_i\ := \$v5583\(0 to 31);
                \$v5587\ := X"0000000" & X"2";
                \$v5585\ := "0000" & \$v5587\;
                \$v5586\ := \$v5585\(0 to 3);
                \$v5584\ := \$v5585\(4 to 35);
                case \$v5586\ is
                when "0000" =>
                  \$13814\ := eclat_false;
                when "0001" =>
                  \$13868_j\ := \$v5584\(0 to 31);
                  \$13814\ := eclat_eq(\$13865_i\ & \$13868_j\);
                when others =>
                  
                end case;
                \$v5582\ := \$13814\;
                if \$v5582\(0) = '1' then
                  \$v5574\ := \$$10700_pc_ptr_take\;
                  if \$v5574\(0) = '1' then
                    state_var7021 <= q_wait5573;
                  else
                    \$$10700_pc_ptr_take\(0) := '1';
                    \$$10700_pc_ptr\ <= 0;
                    state_var7021 <= pause_getI5571;
                  end if;
                else
                  \$v5580\ := \$10793\(36 to 71);
                  \$v5581\ := \$v5580\(0 to 3);
                  \$v5579\ := \$v5580\(4 to 35);
                  case \$v5581\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't int_of_triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$13821_forever3163281\;
                  when "0000" =>
                    \$13829_i\ := \$v5579\(0 to 31);
                    \$13816\ := \$13829_i\;
                    \$v5578\ := \$$10700_pc_ptr_take\;
                    if \$v5578\(0) = '1' then
                      state_var7021 <= q_wait5577;
                    else
                      \$$10700_pc_ptr_take\(0) := '1';
                      \$$10700_pc_ptr_write\ <= 0;
                      \$$10700_pc_write_request\ <= '1';
                      \$$10700_pc_write\ <= \$13816\;
                      state_var7021 <= pause_setI5575;
                    end if;
                  when others =>
                    
                  end case;
                end if;
              when "0000" =>
                \$13869_i\ := \$v5583\(0 to 31);
                \$v5591\ := X"0000000" & X"2";
                \$v5589\ := "0000" & \$v5591\;
                \$v5590\ := \$v5589\(0 to 3);
                \$v5588\ := \$v5589\(4 to 35);
                case \$v5590\ is
                when "0001" =>
                  \$13814\ := eclat_false;
                when "0000" =>
                  \$13872_j\ := \$v5588\(0 to 31);
                  \$13814\ := eclat_eq(\$13869_i\ & \$13872_j\);
                when others =>
                  
                end case;
                \$v5582\ := \$13814\;
                if \$v5582\(0) = '1' then
                  \$v5574\ := \$$10700_pc_ptr_take\;
                  if \$v5574\(0) = '1' then
                    state_var7021 <= q_wait5573;
                  else
                    \$$10700_pc_ptr_take\(0) := '1';
                    \$$10700_pc_ptr\ <= 0;
                    state_var7021 <= pause_getI5571;
                  end if;
                else
                  \$v5580\ := \$10793\(36 to 71);
                  \$v5581\ := \$v5580\(0 to 3);
                  \$v5579\ := \$v5580\(4 to 35);
                  case \$v5581\ is
                  when "0001" =>
                    eclat_print_string(of_string("Fatal error : "));
                    
                    eclat_print_string(of_string("can't int_of_triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var7021 <= \$13821_forever3163281\;
                  when "0000" =>
                    \$13829_i\ := \$v5579\(0 to 31);
                    \$13816\ := \$13829_i\;
                    \$v5578\ := \$$10700_pc_ptr_take\;
                    if \$v5578\(0) = '1' then
                      state_var7021 <= q_wait5577;
                    else
                      \$$10700_pc_ptr_take\(0) := '1';
                      \$$10700_pc_ptr_write\ <= 0;
                      \$$10700_pc_write_request\ <= '1';
                      \$$10700_pc_write\ <= \$13816\;
                      state_var7021 <= pause_setI5575;
                    end if;
                  when others =>
                    
                  end case;
                end if;
              when others =>
                
              end case;
            when pause_setII5624 =>
              \$$10697_stack_ptr_take\(0) := '0';
              state_var7021 <= \$10778_run286\;
            when pause_setII5630 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5626\ := \$$10697_stack_ptr_take\;
              if \$v5626\(0) = '1' then
                state_var7021 <= q_wait5625;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$10767_j\;
                state_var7021 <= pause_setI5623;
              end if;
            when pause_setII5637 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5632\ := \$$10696_ram_ptr_take\;
              if \$v5632\(0) = '1' then
                state_var7021 <= q_wait5631;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5627\ := X"0000000" & X"0";
                \$v5628\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10767_j\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5627\ & "0001" & \$v5628\ & "0000" & \$10763_i\;
                state_var7021 <= pause_setI5629;
              end if;
            when pause_setII5649 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5647\ := \$$10702_brk_ptr_take\;
              if \$v5647\(0) = '1' then
                state_var7021 <= q_wait5646;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5644;
              end if;
            when pause_setII5674 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5672\ := \$$10702_brk_ptr_take\;
              if \$v5672\(0) = '1' then
                state_var7021 <= q_wait5671;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5669;
              end if;
            when pause_setII5691 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v5689\ := \$$10702_brk_ptr_take\;
              if \$v5689\(0) = '1' then
                state_var7021 <= q_wait5688;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5686;
              end if;
            when pause_setII5711 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5707\ := \$$10699_symtbl_ptr_take\;
              if \$v5707\(0) = '1' then
                state_var7021 <= q_wait5706;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5704;
              end if;
            when pause_setII5742 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v5740\ := \$$10699_symtbl_ptr_take\;
              if \$v5740\(0) = '1' then
                state_var7021 <= q_wait5739;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5737;
              end if;
            when pause_setII5762 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5758\ := \$$10699_symtbl_ptr_take\;
              if \$v5758\(0) = '1' then
                state_var7021 <= q_wait5757;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5755;
              end if;
            when pause_setII5793 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v5791\ := \$$10699_symtbl_ptr_take\;
              if \$v5791\(0) = '1' then
                state_var7021 <= q_wait5790;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5788;
              end if;
            when pause_setII5813 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5809\ := \$$10699_symtbl_ptr_take\;
              if \$v5809\(0) = '1' then
                state_var7021 <= q_wait5808;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5806;
              end if;
            when pause_setII5844 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v5842\ := \$$10699_symtbl_ptr_take\;
              if \$v5842\(0) = '1' then
                state_var7021 <= q_wait5841;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5839;
              end if;
            when pause_setII5863 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5860\ := \$$10699_symtbl_ptr_take\;
              if \$v5860\(0) = '1' then
                state_var7021 <= q_wait5859;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5857;
              end if;
            when pause_setII5900 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5896\ := \$$10698_heap_ptr_take\;
              if \$v5896\(0) = '1' then
                state_var7021 <= q_wait5895;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5893;
              end if;
            when pause_setII5908 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v5906\ := \$$10698_heap_ptr_take\;
              if \$v5906\(0) = '1' then
                state_var7021 <= q_wait5905;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5903;
              end if;
            when pause_setII5920 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v5918\ := \$$10702_brk_ptr_take\;
              if \$v5918\(0) = '1' then
                state_var7021 <= q_wait5917;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5915;
              end if;
            when pause_setII5941 =>
              \$$10700_pc_ptr_take\(0) := '0';
              \$v5939\ := \$$10699_symtbl_ptr_take\;
              if \$v5939\(0) = '1' then
                state_var7021 <= q_wait5938;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5936;
              end if;
            when pause_setII5967 =>
              \$$10696_ram_ptr_take\(0) := '0';
              state_var7021 <= \$14481_decode_loop310\;
            when pause_setII5992 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v5989\ := \$$10698_heap_ptr_take\;
              if \$v5989\(0) = '1' then
                state_var7021 <= q_wait5988;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5986;
              end if;
            when pause_setII6000 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v5998\ := \$$10698_heap_ptr_take\;
              if \$v5998\(0) = '1' then
                state_var7021 <= q_wait5997;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5995;
              end if;
            when pause_setII6012 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6010\ := \$$10702_brk_ptr_take\;
              if \$v6010\(0) = '1' then
                state_var7021 <= q_wait6009;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6007;
              end if;
            when pause_setII6040 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$15068_opnd\ := \$15063\(0 to 35);
              \$v6038\ := \$$10697_stack_ptr_take\;
              if \$v6038\(0) = '1' then
                state_var7021 <= q_wait6037;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6035;
              end if;
            when pause_setII6056 =>
              \$$10696_ram_ptr_take\(0) := '0';
              state_var7021 <= \$14481_decode_loop310\;
            when pause_setII6081 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6078\ := \$$10698_heap_ptr_take\;
              if \$v6078\(0) = '1' then
                state_var7021 <= q_wait6077;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6075;
              end if;
            when pause_setII6089 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v6087\ := \$$10698_heap_ptr_take\;
              if \$v6087\(0) = '1' then
                state_var7021 <= q_wait6086;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6084;
              end if;
            when pause_setII6101 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6099\ := \$$10702_brk_ptr_take\;
              if \$v6099\(0) = '1' then
                state_var7021 <= q_wait6098;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6096;
              end if;
            when pause_setII6143 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6139\ := \$$10698_heap_ptr_take\;
              if \$v6139\(0) = '1' then
                state_var7021 <= q_wait6138;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6136;
              end if;
            when pause_setII6151 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v6149\ := \$$10698_heap_ptr_take\;
              if \$v6149\(0) = '1' then
                state_var7021 <= q_wait6148;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6146;
              end if;
            when pause_setII6163 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6161\ := \$$10702_brk_ptr_take\;
              if \$v6161\(0) = '1' then
                state_var7021 <= q_wait6160;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6158;
              end if;
            when pause_setII6185 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6182\ := \$$10698_heap_ptr_take\;
              if \$v6182\(0) = '1' then
                state_var7021 <= q_wait6181;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6179;
              end if;
            when pause_setII6193 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v6191\ := \$$10698_heap_ptr_take\;
              if \$v6191\(0) = '1' then
                state_var7021 <= q_wait6190;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6188;
              end if;
            when pause_setII6205 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6203\ := \$$10702_brk_ptr_take\;
              if \$v6203\(0) = '1' then
                state_var7021 <= q_wait6202;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6200;
              end if;
            when pause_setII6222 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$14648_ty\ := \$14643\(0 to 35);
              \$v6220\ := \$$10702_brk_ptr_take\;
              if \$v6220\(0) = '1' then
                state_var7021 <= q_wait6219;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6217;
              end if;
            when pause_setII6238 =>
              \$$10696_ram_ptr_take\(0) := '0';
              state_var7021 <= \$14481_decode_loop310\;
            when pause_setII6263 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6260\ := \$$10698_heap_ptr_take\;
              if \$v6260\(0) = '1' then
                state_var7021 <= q_wait6259;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6257;
              end if;
            when pause_setII6271 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v6269\ := \$$10698_heap_ptr_take\;
              if \$v6269\(0) = '1' then
                state_var7021 <= q_wait6268;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6266;
              end if;
            when pause_setII6283 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6281\ := \$$10702_brk_ptr_take\;
              if \$v6281\(0) = '1' then
                state_var7021 <= q_wait6280;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6278;
              end if;
            when pause_setII6334 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14949_x\ := eclat_if(eclat_lt(eclat_sub(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$14947\,32) & X"000000" & X"23") & X"0000000" & X"0") & X"000000" & X"39" & eclat_sub(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$14947\,32) & X"000000" & X"23"));
              \$v6332\ := eclat_lt(\$14949_x\ & X"000000" & X"2e");
              if \$v6332\(0) = '1' then
                \$14939_get_int268_result\ := eclat_add(\$14949_x\ & eclat_mult(\$14939_get_int268_arg\(0 to 31) & X"000000" & X"2e"));
                \$14936\ := \$14939_get_int268_result\;
                \$14533_opnd\ := "0001" & \$14936\;
                \$v6310\ := eclat_lt(X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31));
                if \$v6310\(0) = '1' then
                  \$v6235\ := \$$10697_stack_ptr_take\;
                  if \$v6235\(0) = '1' then
                    state_var7021 <= q_wait6234;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI6232;
                  end if;
                else
                  \$v6309\ := \$$10697_stack_ptr_take\;
                  if \$v6309\(0) = '1' then
                    state_var7021 <= q_wait6308;
                  else
                    \$$10697_stack_ptr_take\(0) := '1';
                    \$$10697_stack_ptr\ <= 0;
                    state_var7021 <= pause_getI6306;
                  end if;
                end if;
              else
                \$14939_get_int268_arg\ := eclat_sub(eclat_add(eclat_mult(\$14939_get_int268_arg\(0 to 31) & X"000000" & X"2e") & \$14949_x\) & X"000000" & X"2e") & eclat_unit;
                state_var7021 <= \$14939_get_int268\;
              end if;
            when pause_setII6366 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14913_x\ := eclat_if(eclat_lt(eclat_sub(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$14911\,32) & X"000000" & X"23") & X"0000000" & X"0") & X"000000" & X"39" & eclat_sub(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$14911\,32) & X"000000" & X"23"));
              \$v6364\ := eclat_lt(\$14913_x\ & X"000000" & X"2e");
              if \$v6364\(0) = '1' then
                \$14897_get_int268_result\ := eclat_add(\$14913_x\ & eclat_mult(\$14897_get_int268_arg\(0 to 31) & X"000000" & X"2e"));
                \$14837\ := \$14897_get_int268_result\;
                \$v6363\ := \$$10699_symtbl_ptr_take\;
                if \$v6363\(0) = '1' then
                  state_var7021 <= q_wait6362;
                else
                  \$$10699_symtbl_ptr_take\(0) := '1';
                  \$$10699_symtbl_ptr\ <= 0;
                  state_var7021 <= pause_getI6360;
                end if;
              else
                \$14897_get_int268_arg\ := eclat_sub(eclat_add(eclat_mult(\$14897_get_int268_arg\(0 to 31) & X"000000" & X"2e") & \$14913_x\) & X"000000" & X"2e") & eclat_unit;
                state_var7021 <= \$14897_get_int268\;
              end if;
            when pause_setII6382 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6378\ := eclat_lt(\$14511_loop311_arg\(32 to 63) & eclat_vector_get(X"000000" & X"14" & X"000000" & X"1e" & X"0000000" & X"0" & X"0000000" & X"a" & X"0000000" & X"b" & X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31),32));
              if \$v6378\(0) = '1' then
                \$v6331\ := eclat_lt(\$14511_loop311_arg\(0 to 31) & X"0000000" & X"3");
                if \$v6331\(0) = '1' then
                  \$v6329\ := \$$10699_symtbl_ptr_take\;
                  if \$v6329\(0) = '1' then
                    state_var7021 <= q_wait6328;
                  else
                    \$$10699_symtbl_ptr_take\(0) := '1';
                    \$$10699_symtbl_ptr\ <= 0;
                    state_var7021 <= pause_getI6326;
                  end if;
                else
                  \$v6330\ := \$14511_loop311_arg\(32 to 63);
                  \$14533_opnd\ := "0001" & \$v6330\;
                  \$v6310\ := eclat_lt(X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31));
                  if \$v6310\(0) = '1' then
                    \$v6235\ := \$$10697_stack_ptr_take\;
                    if \$v6235\(0) = '1' then
                      state_var7021 <= q_wait6234;
                    else
                      \$$10697_stack_ptr_take\(0) := '1';
                      \$$10697_stack_ptr\ <= 0;
                      state_var7021 <= pause_getI6232;
                    end if;
                  else
                    \$v6309\ := \$$10697_stack_ptr_take\;
                    if \$v6309\(0) = '1' then
                      state_var7021 <= q_wait6308;
                    else
                      \$$10697_stack_ptr_take\(0) := '1';
                      \$$10697_stack_ptr\ <= 0;
                      state_var7021 <= pause_getI6306;
                    end if;
                  end if;
                end if;
              else
                \$v6377\ := eclat_eq(\$14511_loop311_arg\(32 to 63) & eclat_vector_get(X"000000" & X"14" & X"000000" & X"1e" & X"0000000" & X"0" & X"0000000" & X"a" & X"0000000" & X"b" & X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31),32));
                if \$v6377\(0) = '1' then
                  \$14939_get_int268_arg\ := X"0000000" & X"0" & eclat_unit;
                  state_var7021 <= \$14939_get_int268\;
                else
                  \$14897_get_int268_arg\ := eclat_sub(eclat_sub(\$14511_loop311_arg\(32 to 63) & eclat_vector_get(X"000000" & X"14" & X"000000" & X"1e" & X"0000000" & X"0" & X"0000000" & X"a" & X"0000000" & X"b" & X"0000000" & X"4" & \$14511_loop311_arg\(0 to 31),32)) & X"0000000" & X"1") & eclat_unit;
                  state_var7021 <= \$14897_get_int268\;
                end if;
              end if;
            when pause_setII6390 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v6388\ := \$$10697_stack_ptr_take\;
              if \$v6388\(0) = '1' then
                state_var7021 <= q_wait6387;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6385;
              end if;
            when pause_setII6406 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6404\ := \$$10702_brk_ptr_take\;
              if \$v6404\(0) = '1' then
                state_var7021 <= q_wait6403;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6401;
              end if;
            when pause_setII6426 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$14500_x\ := eclat_if(eclat_lt(eclat_sub(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$14498\,32) & X"000000" & X"23") & X"0000000" & X"0") & X"000000" & X"39" & eclat_sub(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$14498\,32) & X"000000" & X"23"));
              \$14511_loop311_arg\ := X"0000000" & X"0" & \$14500_x\ & \$14500_x\ & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var7021 <= \$14511_loop311\;
            when pause_setII6443 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6440\ := \$$10699_symtbl_ptr_take\;
              if \$v6440\(0) = '1' then
                state_var7021 <= q_wait6439;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6437;
              end if;
            when pause_setII6451 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6449\ := \$$10699_symtbl_ptr_take\;
              if \$v6449\(0) = '1' then
                state_var7021 <= q_wait6448;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6446;
              end if;
            when pause_setII6463 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6461\ := \$$10702_brk_ptr_take\;
              if \$v6461\(0) = '1' then
                state_var7021 <= q_wait6460;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6458;
              end if;
            when pause_setII6486 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6482\ := \$$10699_symtbl_ptr_take\;
              if \$v6482\(0) = '1' then
                state_var7021 <= q_wait6481;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6479;
              end if;
            when pause_setII6494 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6492\ := \$$10699_symtbl_ptr_take\;
              if \$v6492\(0) = '1' then
                state_var7021 <= q_wait6491;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6489;
              end if;
            when pause_setII6506 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6504\ := \$$10702_brk_ptr_take\;
              if \$v6504\(0) = '1' then
                state_var7021 <= q_wait6503;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6501;
              end if;
            when pause_setII6529 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6525\ := \$$10699_symtbl_ptr_take\;
              if \$v6525\(0) = '1' then
                state_var7021 <= q_wait6524;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6522;
              end if;
            when pause_setII6537 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6535\ := \$$10699_symtbl_ptr_take\;
              if \$v6535\(0) = '1' then
                state_var7021 <= q_wait6534;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6532;
              end if;
            when pause_setII6549 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6547\ := \$$10702_brk_ptr_take\;
              if \$v6547\(0) = '1' then
                state_var7021 <= q_wait6546;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6544;
              end if;
            when pause_setII6607 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6604\ := \$$10699_symtbl_ptr_take\;
              if \$v6604\(0) = '1' then
                state_var7021 <= q_wait6603;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6601;
              end if;
            when pause_setII6615 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6613\ := \$$10699_symtbl_ptr_take\;
              if \$v6613\(0) = '1' then
                state_var7021 <= q_wait6612;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6610;
              end if;
            when pause_setII6627 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6625\ := \$$10702_brk_ptr_take\;
              if \$v6625\(0) = '1' then
                state_var7021 <= q_wait6624;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6622;
              end if;
            when pause_setII6650 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6646\ := \$$10699_symtbl_ptr_take\;
              if \$v6646\(0) = '1' then
                state_var7021 <= q_wait6645;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6643;
              end if;
            when pause_setII6658 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6656\ := \$$10699_symtbl_ptr_take\;
              if \$v6656\(0) = '1' then
                state_var7021 <= q_wait6655;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6653;
              end if;
            when pause_setII6670 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6668\ := \$$10702_brk_ptr_take\;
              if \$v6668\(0) = '1' then
                state_var7021 <= q_wait6667;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6665;
              end if;
            when pause_setII6692 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6689\ := \$$10699_symtbl_ptr_take\;
              if \$v6689\(0) = '1' then
                state_var7021 <= q_wait6688;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6686;
              end if;
            when pause_setII6700 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6698\ := \$$10699_symtbl_ptr_take\;
              if \$v6698\(0) = '1' then
                state_var7021 <= q_wait6697;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6695;
              end if;
            when pause_setII6712 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6710\ := \$$10702_brk_ptr_take\;
              if \$v6710\(0) = '1' then
                state_var7021 <= q_wait6709;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6707;
              end if;
            when pause_setII6768 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6765\ := \$$10699_symtbl_ptr_take\;
              if \$v6765\(0) = '1' then
                state_var7021 <= q_wait6764;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6762;
              end if;
            when pause_setII6776 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6774\ := \$$10699_symtbl_ptr_take\;
              if \$v6774\(0) = '1' then
                state_var7021 <= q_wait6773;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6771;
              end if;
            when pause_setII6788 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6786\ := \$$10702_brk_ptr_take\;
              if \$v6786\(0) = '1' then
                state_var7021 <= q_wait6785;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6783;
              end if;
            when pause_setII6811 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6807\ := \$$10699_symtbl_ptr_take\;
              if \$v6807\(0) = '1' then
                state_var7021 <= q_wait6806;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6804;
              end if;
            when pause_setII6819 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6817\ := \$$10699_symtbl_ptr_take\;
              if \$v6817\(0) = '1' then
                state_var7021 <= q_wait6816;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6814;
              end if;
            when pause_setII6831 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6829\ := \$$10702_brk_ptr_take\;
              if \$v6829\(0) = '1' then
                state_var7021 <= q_wait6828;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6826;
              end if;
            when pause_setII6853 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6850\ := \$$10699_symtbl_ptr_take\;
              if \$v6850\(0) = '1' then
                state_var7021 <= q_wait6849;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6847;
              end if;
            when pause_setII6861 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v6859\ := \$$10699_symtbl_ptr_take\;
              if \$v6859\(0) = '1' then
                state_var7021 <= q_wait6858;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6856;
              end if;
            when pause_setII6873 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6871\ := \$$10702_brk_ptr_take\;
              if \$v6871\(0) = '1' then
                state_var7021 <= q_wait6870;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6868;
              end if;
            when pause_setII6930 =>
              \$$10696_ram_ptr_take\(0) := '0';
              \$v6926\ := \$$10698_heap_ptr_take\;
              if \$v6926\(0) = '1' then
                state_var7021 <= q_wait6925;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6923;
              end if;
            when pause_setII6938 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v6936\ := \$$10698_heap_ptr_take\;
              if \$v6936\(0) = '1' then
                state_var7021 <= q_wait6935;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6933;
              end if;
            when pause_setII6950 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6948\ := \$$10702_brk_ptr_take\;
              if \$v6948\(0) = '1' then
                state_var7021 <= q_wait6947;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6945;
              end if;
            when pause_setII6969 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$v6967\ := eclat_eq(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$15255\,32) & X"000000" & X"2c");
              if \$v6967\(0) = '1' then
                \$v6761\ := \$$10699_symtbl_ptr_take\;
                if \$v6761\(0) = '1' then
                  state_var7021 <= q_wait6760;
                else
                  \$$10699_symtbl_ptr_take\(0) := '1';
                  \$$10699_symtbl_ptr\ <= 0;
                  state_var7021 <= pause_getI6758;
                end if;
              else
                \$v6966\ := eclat_eq(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$15255\,32) & X"000000" & X"3b");
                if \$v6966\(0) = '1' then
                  \$v6922\ := \$$10699_symtbl_ptr_take\;
                  if \$v6922\(0) = '1' then
                    state_var7021 <= q_wait6921;
                  else
                    \$$10699_symtbl_ptr_take\(0) := '1';
                    \$$10699_symtbl_ptr\ <= 0;
                    state_var7021 <= pause_getI6919;
                  end if;
                else
                  \$v6965\ := \$$10702_brk_ptr_take\;
                  if \$v6965\(0) = '1' then
                    state_var7021 <= q_wait6964;
                  else
                    \$$10702_brk_ptr_take\(0) := '1';
                    \$$10702_brk_ptr\ <= 0;
                    state_var7021 <= pause_getI6962;
                  end if;
                end if;
              end if;
            when pause_setII6984 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$15798_x\ := eclat_if(eclat_lt(eclat_sub(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$15796\,32) & X"000000" & X"23") & X"0000000" & X"0") & X"000000" & X"39" & eclat_sub(eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$15796\,32) & X"000000" & X"23"));
              \$v6982\ := eclat_lt(\$15798_x\ & X"000000" & X"2e");
              if \$v6982\(0) = '1' then
                \$15788_get_int268_result\ := eclat_add(\$15798_x\ & eclat_mult(\$15788_get_int268_arg\(0 to 31) & X"000000" & X"2e"));
                \$10717\ := \$15788_get_int268_result\;
                \$15217_loop1312_arg\ := \$10717\ & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit & eclat_unit;
                state_var7021 <= \$15217_loop1312\;
              else
                \$15788_get_int268_arg\ := eclat_sub(eclat_add(eclat_mult(\$15788_get_int268_arg\(0 to 31) & X"000000" & X"2e") & \$15798_x\) & X"000000" & X"2e") & eclat_unit;
                state_var7021 <= \$15788_get_int268\;
              end if;
            when pause_setII6996 =>
              \$$10695_limit_ptr_take\(0) := '0';
              \$15788_get_int268_arg\ := X"0000000" & X"0" & eclat_unit;
              state_var7021 <= \$15788_get_int268\;
            when pause_setII7000 =>
              \$$10702_brk_ptr_take\(0) := '0';
              \$v6998\ := \$$10695_limit_ptr_take\;
              if \$v6998\(0) = '1' then
                state_var7021 <= q_wait6997;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr_write\ <= 0;
                \$$10695_limit_write_request\ <= '1';
                \$$10695_limit_write\ <= eclat_div(X"0000" & X"2710" & X"0000000" & X"2");
                state_var7021 <= pause_setI6995;
              end if;
            when pause_setII7004 =>
              \$$10701_pos_ptr_take\(0) := '0';
              \$v7002\ := \$$10702_brk_ptr_take\;
              if \$v7002\(0) = '1' then
                state_var7021 <= q_wait7001;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= X"0000000" & X"4";
                state_var7021 <= pause_setI6999;
              end if;
            when pause_setII7008 =>
              \$$10699_symtbl_ptr_take\(0) := '0';
              \$v7006\ := \$$10701_pos_ptr_take\;
              if \$v7006\(0) = '1' then
                state_var7021 <= q_wait7005;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= X"0000000" & X"0";
                state_var7021 <= pause_setI7003;
              end if;
            when pause_setII7012 =>
              \$$10698_heap_ptr_take\(0) := '0';
              \$v7010\ := \$$10699_symtbl_ptr_take\;
              if \$v7010\(0) = '1' then
                state_var7021 <= q_wait7009;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= eclat_sub(X"0000000" & X"0" & X"0000000" & X"1");
                state_var7021 <= pause_setI7007;
              end if;
            when pause_setII7016 =>
              \$$10697_stack_ptr_take\(0) := '0';
              \$v7014\ := \$$10698_heap_ptr_take\;
              if \$v7014\(0) = '1' then
                state_var7021 <= q_wait7013;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= eclat_sub(X"0000000" & X"0" & X"0000000" & X"1");
                state_var7021 <= pause_setI7011;
              end if;
            when q_wait3372 =>
              \$v3373\ := \$$10700_pc_ptr_take\;
              if \$v3373\(0) = '1' then
                state_var7021 <= q_wait3372;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$10853\;
                state_var7021 <= pause_setI3370;
              end if;
            when q_wait3380 =>
              \$v3381\ := \$$10696_ram_ptr_take\;
              if \$v3381\(0) = '1' then
                state_var7021 <= q_wait3380;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$10880_i\));
                state_var7021 <= pause_getI3378;
              end if;
            when q_wait3386 =>
              \$v3387\ := \$$10697_stack_ptr_take\;
              if \$v3387\(0) = '1' then
                state_var7021 <= q_wait3386;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$10842\;
                state_var7021 <= pause_setI3384;
              end if;
            when q_wait3394 =>
              \$v3395\ := \$$10696_ram_ptr_take\;
              if \$v3395\(0) = '1' then
                state_var7021 <= q_wait3394;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11098_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11099\(0 to 35) & \$11100\(36 to 71) & \$10814\(72 to 107);
                state_var7021 <= pause_setI3392;
              end if;
            when q_wait3399 =>
              \$v3400\ := \$$10696_ram_ptr_take\;
              if \$v3400\(0) = '1' then
                state_var7021 <= q_wait3399;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11121_i\));
                state_var7021 <= pause_getI3397;
              end if;
            when q_wait3406 =>
              \$v3407\ := \$$10696_ram_ptr_take\;
              if \$v3407\(0) = '1' then
                state_var7021 <= q_wait3406;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11134_i\));
                state_var7021 <= pause_getI3404;
              end if;
            when q_wait3415 =>
              \$v3416\ := \$$10696_ram_ptr_take\;
              if \$v3416\(0) = '1' then
                state_var7021 <= q_wait3415;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11147_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$11084\ & \$11148\(36 to 71) & \$11149\(72 to 107);
                state_var7021 <= pause_setI3413;
              end if;
            when q_wait3420 =>
              \$v3421\ := \$$10696_ram_ptr_take\;
              if \$v3421\(0) = '1' then
                state_var7021 <= q_wait3420;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11172_i\));
                state_var7021 <= pause_getI3418;
              end if;
            when q_wait3427 =>
              \$v3428\ := \$$10696_ram_ptr_take\;
              if \$v3428\(0) = '1' then
                state_var7021 <= q_wait3427;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11185_i\));
                state_var7021 <= pause_getI3425;
              end if;
            when q_wait3435 =>
              \$v3436\ := \$$10697_stack_ptr_take\;
              if \$v3436\(0) = '1' then
                state_var7021 <= q_wait3435;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3433;
              end if;
            when q_wait3440 =>
              \$v3441\ := \$$10696_ram_ptr_take\;
              if \$v3441\(0) = '1' then
                state_var7021 <= q_wait3440;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10913_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$10914\(0 to 35) & \$10915\(36 to 71) & \$10900\(72 to 107);
                state_var7021 <= pause_setI3438;
              end if;
            when q_wait3445 =>
              \$v3446\ := \$$10696_ram_ptr_take\;
              if \$v3446\(0) = '1' then
                state_var7021 <= q_wait3445;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$10940_i\));
                state_var7021 <= pause_getI3443;
              end if;
            when q_wait3452 =>
              \$v3453\ := \$$10696_ram_ptr_take\;
              if \$v3453\(0) = '1' then
                state_var7021 <= q_wait3452;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$10953_i\));
                state_var7021 <= pause_getI3450;
              end if;
            when q_wait3461 =>
              \$v3462\ := \$$10696_ram_ptr_take\;
              if \$v3462\(0) = '1' then
                state_var7021 <= q_wait3461;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$10966_i\));
                state_var7021 <= pause_getI3459;
              end if;
            when q_wait3468 =>
              \$v3469\ := \$$10696_ram_ptr_take\;
              if \$v3469\(0) = '1' then
                state_var7021 <= q_wait3468;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10979_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$10898\(0 to 35) & \$10980\(36 to 71) & \$10981\(72 to 107);
                state_var7021 <= pause_setI3466;
              end if;
            when q_wait3473 =>
              \$v3474\ := \$$10696_ram_ptr_take\;
              if \$v3474\(0) = '1' then
                state_var7021 <= q_wait3473;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11006_i\));
                state_var7021 <= pause_getI3471;
              end if;
            when q_wait3480 =>
              \$v3481\ := \$$10696_ram_ptr_take\;
              if \$v3481\(0) = '1' then
                state_var7021 <= q_wait3480;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11019_i\));
                state_var7021 <= pause_getI3478;
              end if;
            when q_wait3489 =>
              \$v3490\ := \$$10696_ram_ptr_take\;
              if \$v3490\(0) = '1' then
                state_var7021 <= q_wait3489;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11032_i\));
                state_var7021 <= pause_getI3487;
              end if;
            when q_wait3496 =>
              \$v3497\ := \$$10696_ram_ptr_take\;
              if \$v3497\(0) = '1' then
                state_var7021 <= q_wait3496;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11065_i\));
                state_var7021 <= pause_getI3494;
              end if;
            when q_wait3507 =>
              \$v3508\ := \$$10696_ram_ptr_take\;
              if \$v3508\(0) = '1' then
                state_var7021 <= q_wait3507;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11081_i\));
                state_var7021 <= pause_getI3505;
              end if;
            when q_wait3513 =>
              \$v3514\ := \$$10697_stack_ptr_take\;
              if \$v3514\(0) = '1' then
                state_var7021 <= q_wait3513;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3511;
              end if;
            when q_wait3521 =>
              \$v3522\ := \$$10698_heap_ptr_take\;
              if \$v3522\(0) = '1' then
                state_var7021 <= q_wait3521;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3519;
              end if;
            when q_wait3526 =>
              \$v3527\ := \$$10696_ram_ptr_take\;
              if \$v3527\(0) = '1' then
                state_var7021 <= q_wait3526;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3523\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11230\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11219\ & \$11196_loop2913158_arg\(32 to 67) & "0001" & \$v3523\;
                state_var7021 <= pause_setI3524;
              end if;
            when q_wait3530 =>
              \$v3531\ := \$$10698_heap_ptr_take\;
              if \$v3531\(0) = '1' then
                state_var7021 <= q_wait3530;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3528;
              end if;
            when q_wait3534 =>
              \$v3535\ := \$$10698_heap_ptr_take\;
              if \$v3535\(0) = '1' then
                state_var7021 <= q_wait3534;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11228_i\;
                state_var7021 <= pause_setI3532;
              end if;
            when q_wait3538 =>
              \$v3539\ := \$$10702_brk_ptr_take\;
              if \$v3539\(0) = '1' then
                state_var7021 <= q_wait3538;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3536;
              end if;
            when q_wait3542 =>
              \$v3543\ := \$$10702_brk_ptr_take\;
              if \$v3543\(0) = '1' then
                state_var7021 <= q_wait3542;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3540;
              end if;
            when q_wait3546 =>
              \$v3547\ := \$$10702_brk_ptr_take\;
              if \$v3547\(0) = '1' then
                state_var7021 <= q_wait3546;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11236\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3544;
              end if;
            when q_wait3550 =>
              \$v3551\ := \$$10702_brk_ptr_take\;
              if \$v3551\(0) = '1' then
                state_var7021 <= q_wait3550;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3548;
              end if;
            when q_wait3555 =>
              \$v3556\ := \$$10695_limit_ptr_take\;
              if \$v3556\(0) = '1' then
                state_var7021 <= q_wait3555;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3553;
              end if;
            when q_wait3559 =>
              \$v3560\ := \$$10702_brk_ptr_take\;
              if \$v3560\(0) = '1' then
                state_var7021 <= q_wait3559;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3557;
              end if;
            when q_wait3563 =>
              \$v3564\ := \$$10697_stack_ptr_take\;
              if \$v3564\(0) = '1' then
                state_var7021 <= q_wait3563;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11218\;
                state_var7021 <= pause_setI3561;
              end if;
            when q_wait3570 =>
              \$v3571\ := \$$10696_ram_ptr_take\;
              if \$v3571\(0) = '1' then
                state_var7021 <= q_wait3570;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11213\));
                state_var7021 <= pause_getI3568;
              end if;
            when q_wait3574 =>
              \$v3575\ := \$$10697_stack_ptr_take\;
              if \$v3575\(0) = '1' then
                state_var7021 <= q_wait3574;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3572;
              end if;
            when q_wait3583 =>
              \$v3584\ := \$$10696_ram_ptr_take\;
              if \$v3584\(0) = '1' then
                state_var7021 <= q_wait3583;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11293_i\));
                state_var7021 <= pause_getI3581;
              end if;
            when q_wait3589 =>
              \$v3590\ := \$$10698_heap_ptr_take\;
              if \$v3590\(0) = '1' then
                state_var7021 <= q_wait3589;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3587;
              end if;
            when q_wait3595 =>
              \$v3596\ := \$$10696_ram_ptr_take\;
              if \$v3596\(0) = '1' then
                state_var7021 <= q_wait3595;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3591\ := X"0000000" & X"0";
                \$v3592\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11296\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v3591\ & \$10818_proc\ & "0001" & \$v3592\;
                state_var7021 <= pause_setI3593;
              end if;
            when q_wait3599 =>
              \$v3600\ := \$$10698_heap_ptr_take\;
              if \$v3600\(0) = '1' then
                state_var7021 <= q_wait3599;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3597;
              end if;
            when q_wait3603 =>
              \$v3604\ := \$$10698_heap_ptr_take\;
              if \$v3604\(0) = '1' then
                state_var7021 <= q_wait3603;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11294_i\;
                state_var7021 <= pause_setI3601;
              end if;
            when q_wait3607 =>
              \$v3608\ := \$$10702_brk_ptr_take\;
              if \$v3608\(0) = '1' then
                state_var7021 <= q_wait3607;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3605;
              end if;
            when q_wait3611 =>
              \$v3612\ := \$$10702_brk_ptr_take\;
              if \$v3612\(0) = '1' then
                state_var7021 <= q_wait3611;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3609;
              end if;
            when q_wait3615 =>
              \$v3616\ := \$$10702_brk_ptr_take\;
              if \$v3616\(0) = '1' then
                state_var7021 <= q_wait3615;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11303\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3613;
              end if;
            when q_wait3619 =>
              \$v3620\ := \$$10702_brk_ptr_take\;
              if \$v3620\(0) = '1' then
                state_var7021 <= q_wait3619;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3617;
              end if;
            when q_wait3624 =>
              \$v3625\ := \$$10695_limit_ptr_take\;
              if \$v3625\(0) = '1' then
                state_var7021 <= q_wait3624;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3622;
              end if;
            when q_wait3628 =>
              \$v3629\ := \$$10702_brk_ptr_take\;
              if \$v3629\(0) = '1' then
                state_var7021 <= q_wait3628;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3626;
              end if;
            when q_wait3632 =>
              \$v3633\ := \$$10700_pc_ptr_take\;
              if \$v3633\(0) = '1' then
                state_var7021 <= q_wait3632;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$11491\;
                state_var7021 <= pause_setI3630;
              end if;
            when q_wait3640 =>
              \$v3641\ := \$$10696_ram_ptr_take\;
              if \$v3641\(0) = '1' then
                state_var7021 <= q_wait3640;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11518_i\));
                state_var7021 <= pause_getI3638;
              end if;
            when q_wait3646 =>
              \$v3647\ := \$$10700_pc_ptr_take\;
              if \$v3647\(0) = '1' then
                state_var7021 <= q_wait3646;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI3644;
              end if;
            when q_wait3650 =>
              \$v3651\ := \$$10700_pc_ptr_take\;
              if \$v3651\(0) = '1' then
                state_var7021 <= q_wait3650;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$11338\;
                state_var7021 <= pause_setI3648;
              end if;
            when q_wait3658 =>
              \$v3659\ := \$$10696_ram_ptr_take\;
              if \$v3659\(0) = '1' then
                state_var7021 <= q_wait3658;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11364_i\));
                state_var7021 <= pause_getI3656;
              end if;
            when q_wait3665 =>
              \$v3666\ := \$$10696_ram_ptr_take\;
              if \$v3666\(0) = '1' then
                state_var7021 <= q_wait3665;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11378_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11379\(0 to 35) & \$11331\(0 to 35) & \$11380\(72 to 107);
                state_var7021 <= pause_setI3663;
              end if;
            when q_wait3670 =>
              \$v3671\ := \$$10696_ram_ptr_take\;
              if \$v3671\(0) = '1' then
                state_var7021 <= q_wait3670;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11406_i\));
                state_var7021 <= pause_getI3668;
              end if;
            when q_wait3677 =>
              \$v3678\ := \$$10696_ram_ptr_take\;
              if \$v3678\(0) = '1' then
                state_var7021 <= q_wait3677;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11420_i\));
                state_var7021 <= pause_getI3675;
              end if;
            when q_wait3686 =>
              \$v3687\ := \$$10696_ram_ptr_take\;
              if \$v3687\(0) = '1' then
                state_var7021 <= q_wait3686;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11433_i\));
                state_var7021 <= pause_getI3684;
              end if;
            when q_wait3692 =>
              \$v3693\ := \$$10697_stack_ptr_take\;
              if \$v3693\(0) = '1' then
                state_var7021 <= q_wait3692;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3690;
              end if;
            when q_wait3697 =>
              \$v3698\ := \$$10696_ram_ptr_take\;
              if \$v3698\(0) = '1' then
                state_var7021 <= q_wait3697;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11466_i\));
                state_var7021 <= pause_getI3695;
              end if;
            when q_wait3708 =>
              \$v3709\ := \$$10696_ram_ptr_take\;
              if \$v3709\(0) = '1' then
                state_var7021 <= q_wait3708;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11482_i\));
                state_var7021 <= pause_getI3706;
              end if;
            when q_wait3714 =>
              \$v3715\ := \$$10697_stack_ptr_take\;
              if \$v3715\(0) = '1' then
                state_var7021 <= q_wait3714;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3712;
              end if;
            when q_wait3723 =>
              \$v3724\ := \$$10696_ram_ptr_take\;
              if \$v3724\(0) = '1' then
                state_var7021 <= q_wait3723;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3720\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11571\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11564_r\ & "0000" & \$11569\ & "0001" & \$v3720\;
                state_var7021 <= pause_setI3721;
              end if;
            when q_wait3727 =>
              \$v3728\ := \$$10697_stack_ptr_take\;
              if \$v3728\(0) = '1' then
                state_var7021 <= q_wait3727;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3725;
              end if;
            when q_wait3731 =>
              \$v3732\ := \$$10697_stack_ptr_take\;
              if \$v3732\(0) = '1' then
                state_var7021 <= q_wait3731;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11568_i\;
                state_var7021 <= pause_setI3729;
              end if;
            when q_wait3735 =>
              \$v3736\ := \$$10697_stack_ptr_take\;
              if \$v3736\(0) = '1' then
                state_var7021 <= q_wait3735;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3733;
              end if;
            when q_wait3739 =>
              \$v3740\ := \$$10702_brk_ptr_take\;
              if \$v3740\(0) = '1' then
                state_var7021 <= q_wait3739;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3737;
              end if;
            when q_wait3743 =>
              \$v3744\ := \$$10702_brk_ptr_take\;
              if \$v3744\(0) = '1' then
                state_var7021 <= q_wait3743;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3741;
              end if;
            when q_wait3747 =>
              \$v3748\ := \$$10702_brk_ptr_take\;
              if \$v3748\(0) = '1' then
                state_var7021 <= q_wait3747;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11576\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3745;
              end if;
            when q_wait3751 =>
              \$v3752\ := \$$10702_brk_ptr_take\;
              if \$v3752\(0) = '1' then
                state_var7021 <= q_wait3751;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3749;
              end if;
            when q_wait3756 =>
              \$v3757\ := \$$10695_limit_ptr_take\;
              if \$v3757\(0) = '1' then
                state_var7021 <= q_wait3756;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3754;
              end if;
            when q_wait3760 =>
              \$v3761\ := \$$10702_brk_ptr_take\;
              if \$v3761\(0) = '1' then
                state_var7021 <= q_wait3760;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3758;
              end if;
            when q_wait3764 =>
              \$v3765\ := \$$10698_heap_ptr_take\;
              if \$v3765\(0) = '1' then
                state_var7021 <= q_wait3764;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3762;
              end if;
            when q_wait3768 =>
              \$v3769\ := \$$10696_ram_ptr_take\;
              if \$v3769\(0) = '1' then
                state_var7021 <= q_wait3768;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11562\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11556_z\ & \$11548_y\ & \$11540_x\;
                state_var7021 <= pause_setI3766;
              end if;
            when q_wait3772 =>
              \$v3773\ := \$$10698_heap_ptr_take\;
              if \$v3773\(0) = '1' then
                state_var7021 <= q_wait3772;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI3770;
              end if;
            when q_wait3776 =>
              \$v3777\ := \$$10698_heap_ptr_take\;
              if \$v3777\(0) = '1' then
                state_var7021 <= q_wait3776;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11560_i\;
                state_var7021 <= pause_setI3774;
              end if;
            when q_wait3780 =>
              \$v3781\ := \$$10702_brk_ptr_take\;
              if \$v3781\(0) = '1' then
                state_var7021 <= q_wait3780;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3778;
              end if;
            when q_wait3784 =>
              \$v3785\ := \$$10702_brk_ptr_take\;
              if \$v3785\(0) = '1' then
                state_var7021 <= q_wait3784;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3782;
              end if;
            when q_wait3788 =>
              \$v3789\ := \$$10702_brk_ptr_take\;
              if \$v3789\(0) = '1' then
                state_var7021 <= q_wait3788;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11596\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3786;
              end if;
            when q_wait3792 =>
              \$v3793\ := \$$10702_brk_ptr_take\;
              if \$v3793\(0) = '1' then
                state_var7021 <= q_wait3792;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3790;
              end if;
            when q_wait3797 =>
              \$v3798\ := \$$10695_limit_ptr_take\;
              if \$v3798\(0) = '1' then
                state_var7021 <= q_wait3797;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3795;
              end if;
            when q_wait3801 =>
              \$v3802\ := \$$10702_brk_ptr_take\;
              if \$v3802\(0) = '1' then
                state_var7021 <= q_wait3801;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3799;
              end if;
            when q_wait3805 =>
              \$v3806\ := \$$10697_stack_ptr_take\;
              if \$v3806\(0) = '1' then
                state_var7021 <= q_wait3805;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11555\;
                state_var7021 <= pause_setI3803;
              end if;
            when q_wait3812 =>
              \$v3813\ := \$$10696_ram_ptr_take\;
              if \$v3813\(0) = '1' then
                state_var7021 <= q_wait3812;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11550\));
                state_var7021 <= pause_getI3810;
              end if;
            when q_wait3816 =>
              \$v3817\ := \$$10697_stack_ptr_take\;
              if \$v3817\(0) = '1' then
                state_var7021 <= q_wait3816;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3814;
              end if;
            when q_wait3820 =>
              \$v3821\ := \$$10697_stack_ptr_take\;
              if \$v3821\(0) = '1' then
                state_var7021 <= q_wait3820;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11547\;
                state_var7021 <= pause_setI3818;
              end if;
            when q_wait3827 =>
              \$v3828\ := \$$10696_ram_ptr_take\;
              if \$v3828\(0) = '1' then
                state_var7021 <= q_wait3827;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11542\));
                state_var7021 <= pause_getI3825;
              end if;
            when q_wait3831 =>
              \$v3832\ := \$$10697_stack_ptr_take\;
              if \$v3832\(0) = '1' then
                state_var7021 <= q_wait3831;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3829;
              end if;
            when q_wait3835 =>
              \$v3836\ := \$$10697_stack_ptr_take\;
              if \$v3836\(0) = '1' then
                state_var7021 <= q_wait3835;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11539\;
                state_var7021 <= pause_setI3833;
              end if;
            when q_wait3842 =>
              \$v3843\ := \$$10696_ram_ptr_take\;
              if \$v3843\(0) = '1' then
                state_var7021 <= q_wait3842;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11534\));
                state_var7021 <= pause_getI3840;
              end if;
            when q_wait3846 =>
              \$v3847\ := \$$10697_stack_ptr_take\;
              if \$v3847\(0) = '1' then
                state_var7021 <= q_wait3846;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3844;
              end if;
            when q_wait3851 =>
              \$v3852\ := \$$10696_ram_ptr_take\;
              if \$v3852\(0) = '1' then
                state_var7021 <= q_wait3851;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3848\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11670\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11663\ & "0000" & \$11668\ & "0001" & \$v3848\;
                state_var7021 <= pause_setI3849;
              end if;
            when q_wait3855 =>
              \$v3856\ := \$$10697_stack_ptr_take\;
              if \$v3856\(0) = '1' then
                state_var7021 <= q_wait3855;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3853;
              end if;
            when q_wait3859 =>
              \$v3860\ := \$$10697_stack_ptr_take\;
              if \$v3860\(0) = '1' then
                state_var7021 <= q_wait3859;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11667_i\;
                state_var7021 <= pause_setI3857;
              end if;
            when q_wait3863 =>
              \$v3864\ := \$$10697_stack_ptr_take\;
              if \$v3864\(0) = '1' then
                state_var7021 <= q_wait3863;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3861;
              end if;
            when q_wait3867 =>
              \$v3868\ := \$$10702_brk_ptr_take\;
              if \$v3868\(0) = '1' then
                state_var7021 <= q_wait3867;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3865;
              end if;
            when q_wait3871 =>
              \$v3872\ := \$$10702_brk_ptr_take\;
              if \$v3872\(0) = '1' then
                state_var7021 <= q_wait3871;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3869;
              end if;
            when q_wait3875 =>
              \$v3876\ := \$$10702_brk_ptr_take\;
              if \$v3876\(0) = '1' then
                state_var7021 <= q_wait3875;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11675\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3873;
              end if;
            when q_wait3879 =>
              \$v3880\ := \$$10702_brk_ptr_take\;
              if \$v3880\(0) = '1' then
                state_var7021 <= q_wait3879;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3877;
              end if;
            when q_wait3884 =>
              \$v3885\ := \$$10695_limit_ptr_take\;
              if \$v3885\(0) = '1' then
                state_var7021 <= q_wait3884;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3882;
              end if;
            when q_wait3888 =>
              \$v3889\ := \$$10702_brk_ptr_take\;
              if \$v3889\(0) = '1' then
                state_var7021 <= q_wait3888;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3886;
              end if;
            when q_wait3892 =>
              \$v3893\ := \$$10697_stack_ptr_take\;
              if \$v3893\(0) = '1' then
                state_var7021 <= q_wait3892;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11662\;
                state_var7021 <= pause_setI3890;
              end if;
            when q_wait3899 =>
              \$v3900\ := \$$10696_ram_ptr_take\;
              if \$v3900\(0) = '1' then
                state_var7021 <= q_wait3899;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11657\));
                state_var7021 <= pause_getI3897;
              end if;
            when q_wait3903 =>
              \$v3904\ := \$$10697_stack_ptr_take\;
              if \$v3904\(0) = '1' then
                state_var7021 <= q_wait3903;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3901;
              end if;
            when q_wait3907 =>
              \$v3908\ := \$$10697_stack_ptr_take\;
              if \$v3908\(0) = '1' then
                state_var7021 <= q_wait3907;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11713\;
                state_var7021 <= pause_setI3905;
              end if;
            when q_wait3914 =>
              \$v3915\ := \$$10696_ram_ptr_take\;
              if \$v3915\(0) = '1' then
                state_var7021 <= q_wait3914;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11708\));
                state_var7021 <= pause_getI3912;
              end if;
            when q_wait3918 =>
              \$v3919\ := \$$10697_stack_ptr_take\;
              if \$v3919\(0) = '1' then
                state_var7021 <= q_wait3918;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3916;
              end if;
            when q_wait3923 =>
              \$v3924\ := \$$10696_ram_ptr_take\;
              if \$v3924\(0) = '1' then
                state_var7021 <= q_wait3923;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3920\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11751\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11736_x\ & "0000" & \$11749\ & "0001" & \$v3920\;
                state_var7021 <= pause_setI3921;
              end if;
            when q_wait3927 =>
              \$v3928\ := \$$10697_stack_ptr_take\;
              if \$v3928\(0) = '1' then
                state_var7021 <= q_wait3927;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3925;
              end if;
            when q_wait3931 =>
              \$v3932\ := \$$10697_stack_ptr_take\;
              if \$v3932\(0) = '1' then
                state_var7021 <= q_wait3931;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11748_i\;
                state_var7021 <= pause_setI3929;
              end if;
            when q_wait3935 =>
              \$v3936\ := \$$10697_stack_ptr_take\;
              if \$v3936\(0) = '1' then
                state_var7021 <= q_wait3935;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3933;
              end if;
            when q_wait3939 =>
              \$v3940\ := \$$10702_brk_ptr_take\;
              if \$v3940\(0) = '1' then
                state_var7021 <= q_wait3939;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3937;
              end if;
            when q_wait3943 =>
              \$v3944\ := \$$10702_brk_ptr_take\;
              if \$v3944\(0) = '1' then
                state_var7021 <= q_wait3943;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3941;
              end if;
            when q_wait3947 =>
              \$v3948\ := \$$10702_brk_ptr_take\;
              if \$v3948\(0) = '1' then
                state_var7021 <= q_wait3947;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11756\ & X"0000000" & X"1");
                state_var7021 <= pause_setI3945;
              end if;
            when q_wait3951 =>
              \$v3952\ := \$$10702_brk_ptr_take\;
              if \$v3952\(0) = '1' then
                state_var7021 <= q_wait3951;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3949;
              end if;
            when q_wait3956 =>
              \$v3957\ := \$$10695_limit_ptr_take\;
              if \$v3957\(0) = '1' then
                state_var7021 <= q_wait3956;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI3954;
              end if;
            when q_wait3960 =>
              \$v3961\ := \$$10702_brk_ptr_take\;
              if \$v3961\(0) = '1' then
                state_var7021 <= q_wait3960;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI3958;
              end if;
            when q_wait3964 =>
              \$v3965\ := \$$10697_stack_ptr_take\;
              if \$v3965\(0) = '1' then
                state_var7021 <= q_wait3964;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11743\;
                state_var7021 <= pause_setI3962;
              end if;
            when q_wait3971 =>
              \$v3972\ := \$$10696_ram_ptr_take\;
              if \$v3972\(0) = '1' then
                state_var7021 <= q_wait3971;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11738\));
                state_var7021 <= pause_getI3969;
              end if;
            when q_wait3975 =>
              \$v3976\ := \$$10697_stack_ptr_take\;
              if \$v3976\(0) = '1' then
                state_var7021 <= q_wait3975;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3973;
              end if;
            when q_wait3979 =>
              \$v3980\ := \$$10697_stack_ptr_take\;
              if \$v3980\(0) = '1' then
                state_var7021 <= q_wait3979;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11735\;
                state_var7021 <= pause_setI3977;
              end if;
            when q_wait3986 =>
              \$v3987\ := \$$10696_ram_ptr_take\;
              if \$v3987\(0) = '1' then
                state_var7021 <= q_wait3986;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11730\));
                state_var7021 <= pause_getI3984;
              end if;
            when q_wait3990 =>
              \$v3991\ := \$$10697_stack_ptr_take\;
              if \$v3991\(0) = '1' then
                state_var7021 <= q_wait3990;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3988;
              end if;
            when q_wait3995 =>
              \$v3996\ := \$$10696_ram_ptr_take\;
              if \$v3996\(0) = '1' then
                state_var7021 <= q_wait3995;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v3992\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11821\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11814\ & "0000" & \$11819\ & "0001" & \$v3992\;
                state_var7021 <= pause_setI3993;
              end if;
            when q_wait3999 =>
              \$v4000\ := \$$10697_stack_ptr_take\;
              if \$v4000\(0) = '1' then
                state_var7021 <= q_wait3999;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI3997;
              end if;
            when q_wait4003 =>
              \$v4004\ := \$$10697_stack_ptr_take\;
              if \$v4004\(0) = '1' then
                state_var7021 <= q_wait4003;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11818_i\;
                state_var7021 <= pause_setI4001;
              end if;
            when q_wait4007 =>
              \$v4008\ := \$$10697_stack_ptr_take\;
              if \$v4008\(0) = '1' then
                state_var7021 <= q_wait4007;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4005;
              end if;
            when q_wait4011 =>
              \$v4012\ := \$$10702_brk_ptr_take\;
              if \$v4012\(0) = '1' then
                state_var7021 <= q_wait4011;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4009;
              end if;
            when q_wait4015 =>
              \$v4016\ := \$$10702_brk_ptr_take\;
              if \$v4016\(0) = '1' then
                state_var7021 <= q_wait4015;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4013;
              end if;
            when q_wait4019 =>
              \$v4020\ := \$$10702_brk_ptr_take\;
              if \$v4020\(0) = '1' then
                state_var7021 <= q_wait4019;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11826\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4017;
              end if;
            when q_wait4023 =>
              \$v4024\ := \$$10702_brk_ptr_take\;
              if \$v4024\(0) = '1' then
                state_var7021 <= q_wait4023;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4021;
              end if;
            when q_wait4028 =>
              \$v4029\ := \$$10695_limit_ptr_take\;
              if \$v4029\(0) = '1' then
                state_var7021 <= q_wait4028;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4026;
              end if;
            when q_wait4032 =>
              \$v4033\ := \$$10702_brk_ptr_take\;
              if \$v4033\(0) = '1' then
                state_var7021 <= q_wait4032;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4030;
              end if;
            when q_wait4036 =>
              \$v4037\ := \$$10698_heap_ptr_take\;
              if \$v4037\(0) = '1' then
                state_var7021 <= q_wait4036;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI4034;
              end if;
            when q_wait4041 =>
              \$v4042\ := \$$10696_ram_ptr_take\;
              if \$v4042\(0) = '1' then
                state_var7021 <= q_wait4041;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4038\ := X"0000000" & X"1";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11848\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11810\(0 to 35) & "0000" & \$11812\ & "0001" & \$v4038\;
                state_var7021 <= pause_setI4039;
              end if;
            when q_wait4045 =>
              \$v4046\ := \$$10698_heap_ptr_take\;
              if \$v4046\(0) = '1' then
                state_var7021 <= q_wait4045;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI4043;
              end if;
            when q_wait4049 =>
              \$v4050\ := \$$10698_heap_ptr_take\;
              if \$v4050\(0) = '1' then
                state_var7021 <= q_wait4049;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$11846_i\;
                state_var7021 <= pause_setI4047;
              end if;
            when q_wait4053 =>
              \$v4054\ := \$$10702_brk_ptr_take\;
              if \$v4054\(0) = '1' then
                state_var7021 <= q_wait4053;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4051;
              end if;
            when q_wait4057 =>
              \$v4058\ := \$$10702_brk_ptr_take\;
              if \$v4058\(0) = '1' then
                state_var7021 <= q_wait4057;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4055;
              end if;
            when q_wait4061 =>
              \$v4062\ := \$$10702_brk_ptr_take\;
              if \$v4062\(0) = '1' then
                state_var7021 <= q_wait4061;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11859\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4059;
              end if;
            when q_wait4065 =>
              \$v4066\ := \$$10702_brk_ptr_take\;
              if \$v4066\(0) = '1' then
                state_var7021 <= q_wait4065;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4063;
              end if;
            when q_wait4070 =>
              \$v4071\ := \$$10695_limit_ptr_take\;
              if \$v4071\(0) = '1' then
                state_var7021 <= q_wait4070;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4068;
              end if;
            when q_wait4074 =>
              \$v4075\ := \$$10702_brk_ptr_take\;
              if \$v4075\(0) = '1' then
                state_var7021 <= q_wait4074;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4072;
              end if;
            when q_wait4078 =>
              \$v4079\ := \$$10697_stack_ptr_take\;
              if \$v4079\(0) = '1' then
                state_var7021 <= q_wait4078;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4076;
              end if;
            when q_wait4083 =>
              \$v4084\ := \$$10696_ram_ptr_take\;
              if \$v4084\(0) = '1' then
                state_var7021 <= q_wait4083;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11889_i\));
                state_var7021 <= pause_getI4081;
              end if;
            when q_wait4089 =>
              \$v4090\ := \$$10697_stack_ptr_take\;
              if \$v4090\(0) = '1' then
                state_var7021 <= q_wait4089;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11808\;
                state_var7021 <= pause_setI4087;
              end if;
            when q_wait4096 =>
              \$v4097\ := \$$10696_ram_ptr_take\;
              if \$v4097\(0) = '1' then
                state_var7021 <= q_wait4096;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11803\));
                state_var7021 <= pause_getI4094;
              end if;
            when q_wait4100 =>
              \$v4101\ := \$$10697_stack_ptr_take\;
              if \$v4101\(0) = '1' then
                state_var7021 <= q_wait4100;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4098;
              end if;
            when q_wait4107 =>
              \$v4108\ := \$$10696_ram_ptr_take\;
              if \$v4108\(0) = '1' then
                state_var7021 <= q_wait4107;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4103\ := X"0000000" & X"1";
                \$v4102\ := X"0000000" & X"2";
                \$v4104\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11919\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= eclat_if(\$11912\ & "0000" & \$v4103\ & "0000" & \$v4102\) & "0000" & \$11917\ & "0001" & \$v4104\;
                state_var7021 <= pause_setI4105;
              end if;
            when q_wait4111 =>
              \$v4112\ := \$$10697_stack_ptr_take\;
              if \$v4112\(0) = '1' then
                state_var7021 <= q_wait4111;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4109;
              end if;
            when q_wait4115 =>
              \$v4116\ := \$$10697_stack_ptr_take\;
              if \$v4116\(0) = '1' then
                state_var7021 <= q_wait4115;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11916_i\;
                state_var7021 <= pause_setI4113;
              end if;
            when q_wait4119 =>
              \$v4120\ := \$$10697_stack_ptr_take\;
              if \$v4120\(0) = '1' then
                state_var7021 <= q_wait4119;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4117;
              end if;
            when q_wait4123 =>
              \$v4124\ := \$$10702_brk_ptr_take\;
              if \$v4124\(0) = '1' then
                state_var7021 <= q_wait4123;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4121;
              end if;
            when q_wait4127 =>
              \$v4128\ := \$$10702_brk_ptr_take\;
              if \$v4128\(0) = '1' then
                state_var7021 <= q_wait4127;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4125;
              end if;
            when q_wait4131 =>
              \$v4132\ := \$$10702_brk_ptr_take\;
              if \$v4132\(0) = '1' then
                state_var7021 <= q_wait4131;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11925\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4129;
              end if;
            when q_wait4135 =>
              \$v4136\ := \$$10702_brk_ptr_take\;
              if \$v4136\(0) = '1' then
                state_var7021 <= q_wait4135;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4133;
              end if;
            when q_wait4140 =>
              \$v4141\ := \$$10695_limit_ptr_take\;
              if \$v4141\(0) = '1' then
                state_var7021 <= q_wait4140;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4138;
              end if;
            when q_wait4144 =>
              \$v4145\ := \$$10702_brk_ptr_take\;
              if \$v4145\(0) = '1' then
                state_var7021 <= q_wait4144;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4142;
              end if;
            when q_wait4151 =>
              \$v4152\ := \$$10697_stack_ptr_take\;
              if \$v4152\(0) = '1' then
                state_var7021 <= q_wait4151;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11910\;
                state_var7021 <= pause_setI4149;
              end if;
            when q_wait4158 =>
              \$v4159\ := \$$10696_ram_ptr_take\;
              if \$v4159\(0) = '1' then
                state_var7021 <= q_wait4158;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11905\));
                state_var7021 <= pause_getI4156;
              end if;
            when q_wait4162 =>
              \$v4163\ := \$$10697_stack_ptr_take\;
              if \$v4163\(0) = '1' then
                state_var7021 <= q_wait4162;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4160;
              end if;
            when q_wait4167 =>
              \$v4168\ := \$$10696_ram_ptr_take\;
              if \$v4168\(0) = '1' then
                state_var7021 <= q_wait4167;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4164\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$11975\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$11968\(0 to 35) & "0000" & \$11973\ & "0001" & \$v4164\;
                state_var7021 <= pause_setI4165;
              end if;
            when q_wait4171 =>
              \$v4172\ := \$$10697_stack_ptr_take\;
              if \$v4172\(0) = '1' then
                state_var7021 <= q_wait4171;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4169;
              end if;
            when q_wait4175 =>
              \$v4176\ := \$$10697_stack_ptr_take\;
              if \$v4176\(0) = '1' then
                state_var7021 <= q_wait4175;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11972_i\;
                state_var7021 <= pause_setI4173;
              end if;
            when q_wait4179 =>
              \$v4180\ := \$$10697_stack_ptr_take\;
              if \$v4180\(0) = '1' then
                state_var7021 <= q_wait4179;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4177;
              end if;
            when q_wait4183 =>
              \$v4184\ := \$$10702_brk_ptr_take\;
              if \$v4184\(0) = '1' then
                state_var7021 <= q_wait4183;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4181;
              end if;
            when q_wait4187 =>
              \$v4188\ := \$$10702_brk_ptr_take\;
              if \$v4188\(0) = '1' then
                state_var7021 <= q_wait4187;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4185;
              end if;
            when q_wait4191 =>
              \$v4192\ := \$$10702_brk_ptr_take\;
              if \$v4192\(0) = '1' then
                state_var7021 <= q_wait4191;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$11984\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4189;
              end if;
            when q_wait4195 =>
              \$v4196\ := \$$10702_brk_ptr_take\;
              if \$v4196\(0) = '1' then
                state_var7021 <= q_wait4195;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4193;
              end if;
            when q_wait4200 =>
              \$v4201\ := \$$10695_limit_ptr_take\;
              if \$v4201\(0) = '1' then
                state_var7021 <= q_wait4200;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4198;
              end if;
            when q_wait4204 =>
              \$v4205\ := \$$10702_brk_ptr_take\;
              if \$v4205\(0) = '1' then
                state_var7021 <= q_wait4204;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4202;
              end if;
            when q_wait4209 =>
              \$v4210\ := \$$10696_ram_ptr_take\;
              if \$v4210\(0) = '1' then
                state_var7021 <= q_wait4209;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12014_i\));
                state_var7021 <= pause_getI4207;
              end if;
            when q_wait4215 =>
              \$v4216\ := \$$10697_stack_ptr_take\;
              if \$v4216\(0) = '1' then
                state_var7021 <= q_wait4215;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$11966\;
                state_var7021 <= pause_setI4213;
              end if;
            when q_wait4222 =>
              \$v4223\ := \$$10696_ram_ptr_take\;
              if \$v4223\(0) = '1' then
                state_var7021 <= q_wait4222;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$11961\));
                state_var7021 <= pause_getI4220;
              end if;
            when q_wait4226 =>
              \$v4227\ := \$$10697_stack_ptr_take\;
              if \$v4227\(0) = '1' then
                state_var7021 <= q_wait4226;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4224;
              end if;
            when q_wait4231 =>
              \$v4232\ := \$$10696_ram_ptr_take\;
              if \$v4232\(0) = '1' then
                state_var7021 <= q_wait4231;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4228\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12044\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12037\(36 to 71) & "0000" & \$12042\ & "0001" & \$v4228\;
                state_var7021 <= pause_setI4229;
              end if;
            when q_wait4235 =>
              \$v4236\ := \$$10697_stack_ptr_take\;
              if \$v4236\(0) = '1' then
                state_var7021 <= q_wait4235;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4233;
              end if;
            when q_wait4239 =>
              \$v4240\ := \$$10697_stack_ptr_take\;
              if \$v4240\(0) = '1' then
                state_var7021 <= q_wait4239;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12041_i\;
                state_var7021 <= pause_setI4237;
              end if;
            when q_wait4243 =>
              \$v4244\ := \$$10697_stack_ptr_take\;
              if \$v4244\(0) = '1' then
                state_var7021 <= q_wait4243;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4241;
              end if;
            when q_wait4247 =>
              \$v4248\ := \$$10702_brk_ptr_take\;
              if \$v4248\(0) = '1' then
                state_var7021 <= q_wait4247;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4245;
              end if;
            when q_wait4251 =>
              \$v4252\ := \$$10702_brk_ptr_take\;
              if \$v4252\(0) = '1' then
                state_var7021 <= q_wait4251;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4249;
              end if;
            when q_wait4255 =>
              \$v4256\ := \$$10702_brk_ptr_take\;
              if \$v4256\(0) = '1' then
                state_var7021 <= q_wait4255;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12053\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4253;
              end if;
            when q_wait4259 =>
              \$v4260\ := \$$10702_brk_ptr_take\;
              if \$v4260\(0) = '1' then
                state_var7021 <= q_wait4259;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4257;
              end if;
            when q_wait4264 =>
              \$v4265\ := \$$10695_limit_ptr_take\;
              if \$v4265\(0) = '1' then
                state_var7021 <= q_wait4264;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4262;
              end if;
            when q_wait4268 =>
              \$v4269\ := \$$10702_brk_ptr_take\;
              if \$v4269\(0) = '1' then
                state_var7021 <= q_wait4268;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4266;
              end if;
            when q_wait4273 =>
              \$v4274\ := \$$10696_ram_ptr_take\;
              if \$v4274\(0) = '1' then
                state_var7021 <= q_wait4273;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12083_i\));
                state_var7021 <= pause_getI4271;
              end if;
            when q_wait4279 =>
              \$v4280\ := \$$10697_stack_ptr_take\;
              if \$v4280\(0) = '1' then
                state_var7021 <= q_wait4279;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12035\;
                state_var7021 <= pause_setI4277;
              end if;
            when q_wait4286 =>
              \$v4287\ := \$$10696_ram_ptr_take\;
              if \$v4287\(0) = '1' then
                state_var7021 <= q_wait4286;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12030\));
                state_var7021 <= pause_getI4284;
              end if;
            when q_wait4290 =>
              \$v4291\ := \$$10697_stack_ptr_take\;
              if \$v4291\(0) = '1' then
                state_var7021 <= q_wait4290;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4288;
              end if;
            when q_wait4295 =>
              \$v4296\ := \$$10696_ram_ptr_take\;
              if \$v4296\(0) = '1' then
                state_var7021 <= q_wait4295;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4292\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12113\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12106\(72 to 107) & "0000" & \$12111\ & "0001" & \$v4292\;
                state_var7021 <= pause_setI4293;
              end if;
            when q_wait4299 =>
              \$v4300\ := \$$10697_stack_ptr_take\;
              if \$v4300\(0) = '1' then
                state_var7021 <= q_wait4299;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4297;
              end if;
            when q_wait4303 =>
              \$v4304\ := \$$10697_stack_ptr_take\;
              if \$v4304\(0) = '1' then
                state_var7021 <= q_wait4303;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12110_i\;
                state_var7021 <= pause_setI4301;
              end if;
            when q_wait4307 =>
              \$v4308\ := \$$10697_stack_ptr_take\;
              if \$v4308\(0) = '1' then
                state_var7021 <= q_wait4307;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4305;
              end if;
            when q_wait4311 =>
              \$v4312\ := \$$10702_brk_ptr_take\;
              if \$v4312\(0) = '1' then
                state_var7021 <= q_wait4311;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4309;
              end if;
            when q_wait4315 =>
              \$v4316\ := \$$10702_brk_ptr_take\;
              if \$v4316\(0) = '1' then
                state_var7021 <= q_wait4315;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4313;
              end if;
            when q_wait4319 =>
              \$v4320\ := \$$10702_brk_ptr_take\;
              if \$v4320\(0) = '1' then
                state_var7021 <= q_wait4319;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12122\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4317;
              end if;
            when q_wait4323 =>
              \$v4324\ := \$$10702_brk_ptr_take\;
              if \$v4324\(0) = '1' then
                state_var7021 <= q_wait4323;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4321;
              end if;
            when q_wait4328 =>
              \$v4329\ := \$$10695_limit_ptr_take\;
              if \$v4329\(0) = '1' then
                state_var7021 <= q_wait4328;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4326;
              end if;
            when q_wait4332 =>
              \$v4333\ := \$$10702_brk_ptr_take\;
              if \$v4333\(0) = '1' then
                state_var7021 <= q_wait4332;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4330;
              end if;
            when q_wait4337 =>
              \$v4338\ := \$$10696_ram_ptr_take\;
              if \$v4338\(0) = '1' then
                state_var7021 <= q_wait4337;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12152_i\));
                state_var7021 <= pause_getI4335;
              end if;
            when q_wait4343 =>
              \$v4344\ := \$$10697_stack_ptr_take\;
              if \$v4344\(0) = '1' then
                state_var7021 <= q_wait4343;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12104\;
                state_var7021 <= pause_setI4341;
              end if;
            when q_wait4350 =>
              \$v4351\ := \$$10696_ram_ptr_take\;
              if \$v4351\(0) = '1' then
                state_var7021 <= q_wait4350;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12099\));
                state_var7021 <= pause_getI4348;
              end if;
            when q_wait4354 =>
              \$v4355\ := \$$10697_stack_ptr_take\;
              if \$v4355\(0) = '1' then
                state_var7021 <= q_wait4354;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4352;
              end if;
            when q_wait4359 =>
              \$v4360\ := \$$10696_ram_ptr_take\;
              if \$v4360\(0) = '1' then
                state_var7021 <= q_wait4359;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4356\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12190\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12174_x\ & "0000" & \$12188\ & "0001" & \$v4356\;
                state_var7021 <= pause_setI4357;
              end if;
            when q_wait4363 =>
              \$v4364\ := \$$10697_stack_ptr_take\;
              if \$v4364\(0) = '1' then
                state_var7021 <= q_wait4363;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4361;
              end if;
            when q_wait4367 =>
              \$v4368\ := \$$10697_stack_ptr_take\;
              if \$v4368\(0) = '1' then
                state_var7021 <= q_wait4367;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12187_i\;
                state_var7021 <= pause_setI4365;
              end if;
            when q_wait4371 =>
              \$v4372\ := \$$10697_stack_ptr_take\;
              if \$v4372\(0) = '1' then
                state_var7021 <= q_wait4371;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4369;
              end if;
            when q_wait4375 =>
              \$v4376\ := \$$10702_brk_ptr_take\;
              if \$v4376\(0) = '1' then
                state_var7021 <= q_wait4375;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4373;
              end if;
            when q_wait4379 =>
              \$v4380\ := \$$10702_brk_ptr_take\;
              if \$v4380\(0) = '1' then
                state_var7021 <= q_wait4379;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4377;
              end if;
            when q_wait4383 =>
              \$v4384\ := \$$10702_brk_ptr_take\;
              if \$v4384\(0) = '1' then
                state_var7021 <= q_wait4383;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12195\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4381;
              end if;
            when q_wait4387 =>
              \$v4388\ := \$$10702_brk_ptr_take\;
              if \$v4388\(0) = '1' then
                state_var7021 <= q_wait4387;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4385;
              end if;
            when q_wait4392 =>
              \$v4393\ := \$$10695_limit_ptr_take\;
              if \$v4393\(0) = '1' then
                state_var7021 <= q_wait4392;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4390;
              end if;
            when q_wait4396 =>
              \$v4397\ := \$$10702_brk_ptr_take\;
              if \$v4397\(0) = '1' then
                state_var7021 <= q_wait4396;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4394;
              end if;
            when q_wait4401 =>
              \$v4402\ := \$$10696_ram_ptr_take\;
              if \$v4402\(0) = '1' then
                state_var7021 <= q_wait4401;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12225_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12174_x\ & \$12226\(36 to 71) & \$12227\(72 to 107);
                state_var7021 <= pause_setI4399;
              end if;
            when q_wait4406 =>
              \$v4407\ := \$$10696_ram_ptr_take\;
              if \$v4407\(0) = '1' then
                state_var7021 <= q_wait4406;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12248_i\));
                state_var7021 <= pause_getI4404;
              end if;
            when q_wait4413 =>
              \$v4414\ := \$$10696_ram_ptr_take\;
              if \$v4414\(0) = '1' then
                state_var7021 <= q_wait4413;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12261_i\));
                state_var7021 <= pause_getI4411;
              end if;
            when q_wait4421 =>
              \$v4422\ := \$$10697_stack_ptr_take\;
              if \$v4422\(0) = '1' then
                state_var7021 <= q_wait4421;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12181\;
                state_var7021 <= pause_setI4419;
              end if;
            when q_wait4428 =>
              \$v4429\ := \$$10696_ram_ptr_take\;
              if \$v4429\(0) = '1' then
                state_var7021 <= q_wait4428;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12176\));
                state_var7021 <= pause_getI4426;
              end if;
            when q_wait4432 =>
              \$v4433\ := \$$10697_stack_ptr_take\;
              if \$v4433\(0) = '1' then
                state_var7021 <= q_wait4432;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4430;
              end if;
            when q_wait4436 =>
              \$v4437\ := \$$10697_stack_ptr_take\;
              if \$v4437\(0) = '1' then
                state_var7021 <= q_wait4436;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12173\;
                state_var7021 <= pause_setI4434;
              end if;
            when q_wait4443 =>
              \$v4444\ := \$$10696_ram_ptr_take\;
              if \$v4444\(0) = '1' then
                state_var7021 <= q_wait4443;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12168\));
                state_var7021 <= pause_getI4441;
              end if;
            when q_wait4447 =>
              \$v4448\ := \$$10697_stack_ptr_take\;
              if \$v4448\(0) = '1' then
                state_var7021 <= q_wait4447;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4445;
              end if;
            when q_wait4452 =>
              \$v4453\ := \$$10696_ram_ptr_take\;
              if \$v4453\(0) = '1' then
                state_var7021 <= q_wait4452;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4449\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12313\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12297_x\ & "0000" & \$12311\ & "0001" & \$v4449\;
                state_var7021 <= pause_setI4450;
              end if;
            when q_wait4456 =>
              \$v4457\ := \$$10697_stack_ptr_take\;
              if \$v4457\(0) = '1' then
                state_var7021 <= q_wait4456;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4454;
              end if;
            when q_wait4460 =>
              \$v4461\ := \$$10697_stack_ptr_take\;
              if \$v4461\(0) = '1' then
                state_var7021 <= q_wait4460;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12310_i\;
                state_var7021 <= pause_setI4458;
              end if;
            when q_wait4464 =>
              \$v4465\ := \$$10697_stack_ptr_take\;
              if \$v4465\(0) = '1' then
                state_var7021 <= q_wait4464;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4462;
              end if;
            when q_wait4468 =>
              \$v4469\ := \$$10702_brk_ptr_take\;
              if \$v4469\(0) = '1' then
                state_var7021 <= q_wait4468;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4466;
              end if;
            when q_wait4472 =>
              \$v4473\ := \$$10702_brk_ptr_take\;
              if \$v4473\(0) = '1' then
                state_var7021 <= q_wait4472;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4470;
              end if;
            when q_wait4476 =>
              \$v4477\ := \$$10702_brk_ptr_take\;
              if \$v4477\(0) = '1' then
                state_var7021 <= q_wait4476;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12318\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4474;
              end if;
            when q_wait4480 =>
              \$v4481\ := \$$10702_brk_ptr_take\;
              if \$v4481\(0) = '1' then
                state_var7021 <= q_wait4480;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4478;
              end if;
            when q_wait4485 =>
              \$v4486\ := \$$10695_limit_ptr_take\;
              if \$v4486\(0) = '1' then
                state_var7021 <= q_wait4485;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4483;
              end if;
            when q_wait4489 =>
              \$v4490\ := \$$10702_brk_ptr_take\;
              if \$v4490\(0) = '1' then
                state_var7021 <= q_wait4489;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4487;
              end if;
            when q_wait4494 =>
              \$v4495\ := \$$10696_ram_ptr_take\;
              if \$v4495\(0) = '1' then
                state_var7021 <= q_wait4494;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12348_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12349\(0 to 35) & \$12297_x\ & \$12350\(72 to 107);
                state_var7021 <= pause_setI4492;
              end if;
            when q_wait4499 =>
              \$v4500\ := \$$10696_ram_ptr_take\;
              if \$v4500\(0) = '1' then
                state_var7021 <= q_wait4499;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12371_i\));
                state_var7021 <= pause_getI4497;
              end if;
            when q_wait4506 =>
              \$v4507\ := \$$10696_ram_ptr_take\;
              if \$v4507\(0) = '1' then
                state_var7021 <= q_wait4506;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12384_i\));
                state_var7021 <= pause_getI4504;
              end if;
            when q_wait4514 =>
              \$v4515\ := \$$10697_stack_ptr_take\;
              if \$v4515\(0) = '1' then
                state_var7021 <= q_wait4514;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12304\;
                state_var7021 <= pause_setI4512;
              end if;
            when q_wait4521 =>
              \$v4522\ := \$$10696_ram_ptr_take\;
              if \$v4522\(0) = '1' then
                state_var7021 <= q_wait4521;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12299\));
                state_var7021 <= pause_getI4519;
              end if;
            when q_wait4525 =>
              \$v4526\ := \$$10697_stack_ptr_take\;
              if \$v4526\(0) = '1' then
                state_var7021 <= q_wait4525;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4523;
              end if;
            when q_wait4529 =>
              \$v4530\ := \$$10697_stack_ptr_take\;
              if \$v4530\(0) = '1' then
                state_var7021 <= q_wait4529;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12296\;
                state_var7021 <= pause_setI4527;
              end if;
            when q_wait4536 =>
              \$v4537\ := \$$10696_ram_ptr_take\;
              if \$v4537\(0) = '1' then
                state_var7021 <= q_wait4536;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12291\));
                state_var7021 <= pause_getI4534;
              end if;
            when q_wait4540 =>
              \$v4541\ := \$$10697_stack_ptr_take\;
              if \$v4541\(0) = '1' then
                state_var7021 <= q_wait4540;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4538;
              end if;
            when q_wait4545 =>
              \$v4546\ := \$$10696_ram_ptr_take\;
              if \$v4546\(0) = '1' then
                state_var7021 <= q_wait4545;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4542\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12436\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12420_x\ & "0000" & \$12434\ & "0001" & \$v4542\;
                state_var7021 <= pause_setI4543;
              end if;
            when q_wait4549 =>
              \$v4550\ := \$$10697_stack_ptr_take\;
              if \$v4550\(0) = '1' then
                state_var7021 <= q_wait4549;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4547;
              end if;
            when q_wait4553 =>
              \$v4554\ := \$$10697_stack_ptr_take\;
              if \$v4554\(0) = '1' then
                state_var7021 <= q_wait4553;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12433_i\;
                state_var7021 <= pause_setI4551;
              end if;
            when q_wait4557 =>
              \$v4558\ := \$$10697_stack_ptr_take\;
              if \$v4558\(0) = '1' then
                state_var7021 <= q_wait4557;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4555;
              end if;
            when q_wait4561 =>
              \$v4562\ := \$$10702_brk_ptr_take\;
              if \$v4562\(0) = '1' then
                state_var7021 <= q_wait4561;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4559;
              end if;
            when q_wait4565 =>
              \$v4566\ := \$$10702_brk_ptr_take\;
              if \$v4566\(0) = '1' then
                state_var7021 <= q_wait4565;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4563;
              end if;
            when q_wait4569 =>
              \$v4570\ := \$$10702_brk_ptr_take\;
              if \$v4570\(0) = '1' then
                state_var7021 <= q_wait4569;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12441\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4567;
              end if;
            when q_wait4573 =>
              \$v4574\ := \$$10702_brk_ptr_take\;
              if \$v4574\(0) = '1' then
                state_var7021 <= q_wait4573;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4571;
              end if;
            when q_wait4578 =>
              \$v4579\ := \$$10695_limit_ptr_take\;
              if \$v4579\(0) = '1' then
                state_var7021 <= q_wait4578;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4576;
              end if;
            when q_wait4582 =>
              \$v4583\ := \$$10702_brk_ptr_take\;
              if \$v4583\(0) = '1' then
                state_var7021 <= q_wait4582;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4580;
              end if;
            when q_wait4587 =>
              \$v4588\ := \$$10696_ram_ptr_take\;
              if \$v4588\(0) = '1' then
                state_var7021 <= q_wait4587;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12471_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12472\(0 to 35) & \$12473\(36 to 71) & \$12420_x\;
                state_var7021 <= pause_setI4585;
              end if;
            when q_wait4592 =>
              \$v4593\ := \$$10696_ram_ptr_take\;
              if \$v4593\(0) = '1' then
                state_var7021 <= q_wait4592;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12494_i\));
                state_var7021 <= pause_getI4590;
              end if;
            when q_wait4599 =>
              \$v4600\ := \$$10696_ram_ptr_take\;
              if \$v4600\(0) = '1' then
                state_var7021 <= q_wait4599;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12507_i\));
                state_var7021 <= pause_getI4597;
              end if;
            when q_wait4607 =>
              \$v4608\ := \$$10697_stack_ptr_take\;
              if \$v4608\(0) = '1' then
                state_var7021 <= q_wait4607;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12427\;
                state_var7021 <= pause_setI4605;
              end if;
            when q_wait4614 =>
              \$v4615\ := \$$10696_ram_ptr_take\;
              if \$v4615\(0) = '1' then
                state_var7021 <= q_wait4614;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12422\));
                state_var7021 <= pause_getI4612;
              end if;
            when q_wait4618 =>
              \$v4619\ := \$$10697_stack_ptr_take\;
              if \$v4619\(0) = '1' then
                state_var7021 <= q_wait4618;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4616;
              end if;
            when q_wait4622 =>
              \$v4623\ := \$$10697_stack_ptr_take\;
              if \$v4623\(0) = '1' then
                state_var7021 <= q_wait4622;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12419\;
                state_var7021 <= pause_setI4620;
              end if;
            when q_wait4629 =>
              \$v4630\ := \$$10696_ram_ptr_take\;
              if \$v4630\(0) = '1' then
                state_var7021 <= q_wait4629;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12414\));
                state_var7021 <= pause_getI4627;
              end if;
            when q_wait4633 =>
              \$v4634\ := \$$10697_stack_ptr_take\;
              if \$v4634\(0) = '1' then
                state_var7021 <= q_wait4633;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4631;
              end if;
            when q_wait4640 =>
              \$v4641\ := \$$10696_ram_ptr_take\;
              if \$v4641\(0) = '1' then
                state_var7021 <= q_wait4640;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4636\ := X"0000000" & X"1";
                \$v4635\ := X"0000000" & X"2";
                \$v4637\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12559\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= eclat_if(\$12552\ & "0000" & \$v4636\ & "0000" & \$v4635\) & "0000" & \$12557\ & "0001" & \$v4637\;
                state_var7021 <= pause_setI4638;
              end if;
            when q_wait4644 =>
              \$v4645\ := \$$10697_stack_ptr_take\;
              if \$v4645\(0) = '1' then
                state_var7021 <= q_wait4644;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4642;
              end if;
            when q_wait4648 =>
              \$v4649\ := \$$10697_stack_ptr_take\;
              if \$v4649\(0) = '1' then
                state_var7021 <= q_wait4648;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12556_i\;
                state_var7021 <= pause_setI4646;
              end if;
            when q_wait4652 =>
              \$v4653\ := \$$10697_stack_ptr_take\;
              if \$v4653\(0) = '1' then
                state_var7021 <= q_wait4652;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4650;
              end if;
            when q_wait4656 =>
              \$v4657\ := \$$10702_brk_ptr_take\;
              if \$v4657\(0) = '1' then
                state_var7021 <= q_wait4656;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4654;
              end if;
            when q_wait4660 =>
              \$v4661\ := \$$10702_brk_ptr_take\;
              if \$v4661\(0) = '1' then
                state_var7021 <= q_wait4660;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4658;
              end if;
            when q_wait4664 =>
              \$v4665\ := \$$10702_brk_ptr_take\;
              if \$v4665\(0) = '1' then
                state_var7021 <= q_wait4664;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12565\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4662;
              end if;
            when q_wait4668 =>
              \$v4669\ := \$$10702_brk_ptr_take\;
              if \$v4669\(0) = '1' then
                state_var7021 <= q_wait4668;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4666;
              end if;
            when q_wait4673 =>
              \$v4674\ := \$$10695_limit_ptr_take\;
              if \$v4674\(0) = '1' then
                state_var7021 <= q_wait4673;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4671;
              end if;
            when q_wait4677 =>
              \$v4678\ := \$$10702_brk_ptr_take\;
              if \$v4678\(0) = '1' then
                state_var7021 <= q_wait4677;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4675;
              end if;
            when q_wait4716 =>
              \$v4717\ := \$$10696_ram_ptr_take\;
              if \$v4717\(0) = '1' then
                state_var7021 <= q_wait4716;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12629_i\));
                state_var7021 <= pause_getI4714;
              end if;
            when q_wait4723 =>
              \$v4724\ := \$$10696_ram_ptr_take\;
              if \$v4724\(0) = '1' then
                state_var7021 <= q_wait4723;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12642_i\));
                state_var7021 <= pause_getI4721;
              end if;
            when q_wait4733 =>
              \$v4734\ := \$$10697_stack_ptr_take\;
              if \$v4734\(0) = '1' then
                state_var7021 <= q_wait4733;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12550\;
                state_var7021 <= pause_setI4731;
              end if;
            when q_wait4740 =>
              \$v4741\ := \$$10696_ram_ptr_take\;
              if \$v4741\(0) = '1' then
                state_var7021 <= q_wait4740;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12545\));
                state_var7021 <= pause_getI4738;
              end if;
            when q_wait4744 =>
              \$v4745\ := \$$10697_stack_ptr_take\;
              if \$v4745\(0) = '1' then
                state_var7021 <= q_wait4744;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4742;
              end if;
            when q_wait4748 =>
              \$v4749\ := \$$10697_stack_ptr_take\;
              if \$v4749\(0) = '1' then
                state_var7021 <= q_wait4748;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12542\;
                state_var7021 <= pause_setI4746;
              end if;
            when q_wait4755 =>
              \$v4756\ := \$$10696_ram_ptr_take\;
              if \$v4756\(0) = '1' then
                state_var7021 <= q_wait4755;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12537\));
                state_var7021 <= pause_getI4753;
              end if;
            when q_wait4759 =>
              \$v4760\ := \$$10697_stack_ptr_take\;
              if \$v4760\(0) = '1' then
                state_var7021 <= q_wait4759;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4757;
              end if;
            when q_wait4764 =>
              \$v4765\ := \$$10696_ram_ptr_take\;
              if \$v4765\(0) = '1' then
                state_var7021 <= q_wait4764;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4761\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12694\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12687\ & "0000" & \$12692\ & "0001" & \$v4761\;
                state_var7021 <= pause_setI4762;
              end if;
            when q_wait4768 =>
              \$v4769\ := \$$10697_stack_ptr_take\;
              if \$v4769\(0) = '1' then
                state_var7021 <= q_wait4768;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4766;
              end if;
            when q_wait4772 =>
              \$v4773\ := \$$10697_stack_ptr_take\;
              if \$v4773\(0) = '1' then
                state_var7021 <= q_wait4772;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12691_i\;
                state_var7021 <= pause_setI4770;
              end if;
            when q_wait4776 =>
              \$v4777\ := \$$10697_stack_ptr_take\;
              if \$v4777\(0) = '1' then
                state_var7021 <= q_wait4776;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4774;
              end if;
            when q_wait4780 =>
              \$v4781\ := \$$10702_brk_ptr_take\;
              if \$v4781\(0) = '1' then
                state_var7021 <= q_wait4780;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4778;
              end if;
            when q_wait4784 =>
              \$v4785\ := \$$10702_brk_ptr_take\;
              if \$v4785\(0) = '1' then
                state_var7021 <= q_wait4784;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4782;
              end if;
            when q_wait4788 =>
              \$v4789\ := \$$10702_brk_ptr_take\;
              if \$v4789\(0) = '1' then
                state_var7021 <= q_wait4788;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12699\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4786;
              end if;
            when q_wait4792 =>
              \$v4793\ := \$$10702_brk_ptr_take\;
              if \$v4793\(0) = '1' then
                state_var7021 <= q_wait4792;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4790;
              end if;
            when q_wait4797 =>
              \$v4798\ := \$$10695_limit_ptr_take\;
              if \$v4798\(0) = '1' then
                state_var7021 <= q_wait4797;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4795;
              end if;
            when q_wait4801 =>
              \$v4802\ := \$$10702_brk_ptr_take\;
              if \$v4802\(0) = '1' then
                state_var7021 <= q_wait4801;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4799;
              end if;
            when q_wait4813 =>
              \$v4814\ := \$$10697_stack_ptr_take\;
              if \$v4814\(0) = '1' then
                state_var7021 <= q_wait4813;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12685\;
                state_var7021 <= pause_setI4811;
              end if;
            when q_wait4820 =>
              \$v4821\ := \$$10696_ram_ptr_take\;
              if \$v4821\(0) = '1' then
                state_var7021 <= q_wait4820;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12680\));
                state_var7021 <= pause_getI4818;
              end if;
            when q_wait4824 =>
              \$v4825\ := \$$10697_stack_ptr_take\;
              if \$v4825\(0) = '1' then
                state_var7021 <= q_wait4824;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4822;
              end if;
            when q_wait4828 =>
              \$v4829\ := \$$10697_stack_ptr_take\;
              if \$v4829\(0) = '1' then
                state_var7021 <= q_wait4828;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12677\;
                state_var7021 <= pause_setI4826;
              end if;
            when q_wait4835 =>
              \$v4836\ := \$$10696_ram_ptr_take\;
              if \$v4836\(0) = '1' then
                state_var7021 <= q_wait4835;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12672\));
                state_var7021 <= pause_getI4833;
              end if;
            when q_wait4839 =>
              \$v4840\ := \$$10697_stack_ptr_take\;
              if \$v4840\(0) = '1' then
                state_var7021 <= q_wait4839;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4837;
              end if;
            when q_wait4844 =>
              \$v4845\ := \$$10696_ram_ptr_take\;
              if \$v4845\(0) = '1' then
                state_var7021 <= q_wait4844;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4841\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12793\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12786\ & "0000" & \$12791\ & "0001" & \$v4841\;
                state_var7021 <= pause_setI4842;
              end if;
            when q_wait4848 =>
              \$v4849\ := \$$10697_stack_ptr_take\;
              if \$v4849\(0) = '1' then
                state_var7021 <= q_wait4848;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4846;
              end if;
            when q_wait4852 =>
              \$v4853\ := \$$10697_stack_ptr_take\;
              if \$v4853\(0) = '1' then
                state_var7021 <= q_wait4852;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12790_i\;
                state_var7021 <= pause_setI4850;
              end if;
            when q_wait4856 =>
              \$v4857\ := \$$10697_stack_ptr_take\;
              if \$v4857\(0) = '1' then
                state_var7021 <= q_wait4856;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4854;
              end if;
            when q_wait4860 =>
              \$v4861\ := \$$10702_brk_ptr_take\;
              if \$v4861\(0) = '1' then
                state_var7021 <= q_wait4860;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4858;
              end if;
            when q_wait4864 =>
              \$v4865\ := \$$10702_brk_ptr_take\;
              if \$v4865\(0) = '1' then
                state_var7021 <= q_wait4864;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4862;
              end if;
            when q_wait4868 =>
              \$v4869\ := \$$10702_brk_ptr_take\;
              if \$v4869\(0) = '1' then
                state_var7021 <= q_wait4868;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12798\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4866;
              end if;
            when q_wait4872 =>
              \$v4873\ := \$$10702_brk_ptr_take\;
              if \$v4873\(0) = '1' then
                state_var7021 <= q_wait4872;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4870;
              end if;
            when q_wait4877 =>
              \$v4878\ := \$$10695_limit_ptr_take\;
              if \$v4878\(0) = '1' then
                state_var7021 <= q_wait4877;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4875;
              end if;
            when q_wait4881 =>
              \$v4882\ := \$$10702_brk_ptr_take\;
              if \$v4882\(0) = '1' then
                state_var7021 <= q_wait4881;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4879;
              end if;
            when q_wait4892 =>
              \$v4893\ := \$$10697_stack_ptr_take\;
              if \$v4893\(0) = '1' then
                state_var7021 <= q_wait4892;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12784\;
                state_var7021 <= pause_setI4890;
              end if;
            when q_wait4899 =>
              \$v4900\ := \$$10696_ram_ptr_take\;
              if \$v4900\(0) = '1' then
                state_var7021 <= q_wait4899;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12779\));
                state_var7021 <= pause_getI4897;
              end if;
            when q_wait4903 =>
              \$v4904\ := \$$10697_stack_ptr_take\;
              if \$v4904\(0) = '1' then
                state_var7021 <= q_wait4903;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4901;
              end if;
            when q_wait4907 =>
              \$v4908\ := \$$10697_stack_ptr_take\;
              if \$v4908\(0) = '1' then
                state_var7021 <= q_wait4907;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12776\;
                state_var7021 <= pause_setI4905;
              end if;
            when q_wait4914 =>
              \$v4915\ := \$$10696_ram_ptr_take\;
              if \$v4915\(0) = '1' then
                state_var7021 <= q_wait4914;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12771\));
                state_var7021 <= pause_getI4912;
              end if;
            when q_wait4918 =>
              \$v4919\ := \$$10697_stack_ptr_take\;
              if \$v4919\(0) = '1' then
                state_var7021 <= q_wait4918;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4916;
              end if;
            when q_wait4923 =>
              \$v4924\ := \$$10696_ram_ptr_take\;
              if \$v4924\(0) = '1' then
                state_var7021 <= q_wait4923;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4920\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12893\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12886\ & "0000" & \$12891\ & "0001" & \$v4920\;
                state_var7021 <= pause_setI4921;
              end if;
            when q_wait4927 =>
              \$v4928\ := \$$10697_stack_ptr_take\;
              if \$v4928\(0) = '1' then
                state_var7021 <= q_wait4927;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4925;
              end if;
            when q_wait4931 =>
              \$v4932\ := \$$10697_stack_ptr_take\;
              if \$v4932\(0) = '1' then
                state_var7021 <= q_wait4931;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12890_i\;
                state_var7021 <= pause_setI4929;
              end if;
            when q_wait4935 =>
              \$v4936\ := \$$10697_stack_ptr_take\;
              if \$v4936\(0) = '1' then
                state_var7021 <= q_wait4935;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4933;
              end if;
            when q_wait4939 =>
              \$v4940\ := \$$10702_brk_ptr_take\;
              if \$v4940\(0) = '1' then
                state_var7021 <= q_wait4939;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4937;
              end if;
            when q_wait4943 =>
              \$v4944\ := \$$10702_brk_ptr_take\;
              if \$v4944\(0) = '1' then
                state_var7021 <= q_wait4943;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4941;
              end if;
            when q_wait4947 =>
              \$v4948\ := \$$10702_brk_ptr_take\;
              if \$v4948\(0) = '1' then
                state_var7021 <= q_wait4947;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12898\ & X"0000000" & X"1");
                state_var7021 <= pause_setI4945;
              end if;
            when q_wait4951 =>
              \$v4952\ := \$$10702_brk_ptr_take\;
              if \$v4952\(0) = '1' then
                state_var7021 <= q_wait4951;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4949;
              end if;
            when q_wait4956 =>
              \$v4957\ := \$$10695_limit_ptr_take\;
              if \$v4957\(0) = '1' then
                state_var7021 <= q_wait4956;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI4954;
              end if;
            when q_wait4960 =>
              \$v4961\ := \$$10702_brk_ptr_take\;
              if \$v4961\(0) = '1' then
                state_var7021 <= q_wait4960;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI4958;
              end if;
            when q_wait4971 =>
              \$v4972\ := \$$10697_stack_ptr_take\;
              if \$v4972\(0) = '1' then
                state_var7021 <= q_wait4971;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12884\;
                state_var7021 <= pause_setI4969;
              end if;
            when q_wait4978 =>
              \$v4979\ := \$$10696_ram_ptr_take\;
              if \$v4979\(0) = '1' then
                state_var7021 <= q_wait4978;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12879\));
                state_var7021 <= pause_getI4976;
              end if;
            when q_wait4982 =>
              \$v4983\ := \$$10697_stack_ptr_take\;
              if \$v4983\(0) = '1' then
                state_var7021 <= q_wait4982;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4980;
              end if;
            when q_wait4986 =>
              \$v4987\ := \$$10697_stack_ptr_take\;
              if \$v4987\(0) = '1' then
                state_var7021 <= q_wait4986;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12876\;
                state_var7021 <= pause_setI4984;
              end if;
            when q_wait4993 =>
              \$v4994\ := \$$10696_ram_ptr_take\;
              if \$v4994\(0) = '1' then
                state_var7021 <= q_wait4993;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12871\));
                state_var7021 <= pause_getI4991;
              end if;
            when q_wait4997 =>
              \$v4998\ := \$$10697_stack_ptr_take\;
              if \$v4998\(0) = '1' then
                state_var7021 <= q_wait4997;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI4995;
              end if;
            when q_wait5002 =>
              \$v5003\ := \$$10696_ram_ptr_take\;
              if \$v5003\(0) = '1' then
                state_var7021 <= q_wait5002;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v4999\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$12993\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$12986\ & "0000" & \$12991\ & "0001" & \$v4999\;
                state_var7021 <= pause_setI5000;
              end if;
            when q_wait5006 =>
              \$v5007\ := \$$10697_stack_ptr_take\;
              if \$v5007\(0) = '1' then
                state_var7021 <= q_wait5006;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5004;
              end if;
            when q_wait5010 =>
              \$v5011\ := \$$10697_stack_ptr_take\;
              if \$v5011\(0) = '1' then
                state_var7021 <= q_wait5010;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12990_i\;
                state_var7021 <= pause_setI5008;
              end if;
            when q_wait5014 =>
              \$v5015\ := \$$10697_stack_ptr_take\;
              if \$v5015\(0) = '1' then
                state_var7021 <= q_wait5014;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5012;
              end if;
            when q_wait5018 =>
              \$v5019\ := \$$10702_brk_ptr_take\;
              if \$v5019\(0) = '1' then
                state_var7021 <= q_wait5018;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5016;
              end if;
            when q_wait5022 =>
              \$v5023\ := \$$10702_brk_ptr_take\;
              if \$v5023\(0) = '1' then
                state_var7021 <= q_wait5022;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5020;
              end if;
            when q_wait5026 =>
              \$v5027\ := \$$10702_brk_ptr_take\;
              if \$v5027\(0) = '1' then
                state_var7021 <= q_wait5026;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$12998\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5024;
              end if;
            when q_wait5030 =>
              \$v5031\ := \$$10702_brk_ptr_take\;
              if \$v5031\(0) = '1' then
                state_var7021 <= q_wait5030;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5028;
              end if;
            when q_wait5035 =>
              \$v5036\ := \$$10695_limit_ptr_take\;
              if \$v5036\(0) = '1' then
                state_var7021 <= q_wait5035;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5033;
              end if;
            when q_wait5039 =>
              \$v5040\ := \$$10702_brk_ptr_take\;
              if \$v5040\(0) = '1' then
                state_var7021 <= q_wait5039;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5037;
              end if;
            when q_wait5050 =>
              \$v5051\ := \$$10697_stack_ptr_take\;
              if \$v5051\(0) = '1' then
                state_var7021 <= q_wait5050;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12984\;
                state_var7021 <= pause_setI5048;
              end if;
            when q_wait5057 =>
              \$v5058\ := \$$10696_ram_ptr_take\;
              if \$v5058\(0) = '1' then
                state_var7021 <= q_wait5057;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12979\));
                state_var7021 <= pause_getI5055;
              end if;
            when q_wait5061 =>
              \$v5062\ := \$$10697_stack_ptr_take\;
              if \$v5062\(0) = '1' then
                state_var7021 <= q_wait5061;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5059;
              end if;
            when q_wait5065 =>
              \$v5066\ := \$$10697_stack_ptr_take\;
              if \$v5066\(0) = '1' then
                state_var7021 <= q_wait5065;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$12976\;
                state_var7021 <= pause_setI5063;
              end if;
            when q_wait5072 =>
              \$v5073\ := \$$10696_ram_ptr_take\;
              if \$v5073\(0) = '1' then
                state_var7021 <= q_wait5072;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$12971\));
                state_var7021 <= pause_getI5070;
              end if;
            when q_wait5076 =>
              \$v5077\ := \$$10697_stack_ptr_take\;
              if \$v5077\(0) = '1' then
                state_var7021 <= q_wait5076;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5074;
              end if;
            when q_wait5081 =>
              \$v5082\ := \$$10696_ram_ptr_take\;
              if \$v5082\(0) = '1' then
                state_var7021 <= q_wait5081;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5078\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13093\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13086\ & "0000" & \$13091\ & "0001" & \$v5078\;
                state_var7021 <= pause_setI5079;
              end if;
            when q_wait5085 =>
              \$v5086\ := \$$10697_stack_ptr_take\;
              if \$v5086\(0) = '1' then
                state_var7021 <= q_wait5085;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5083;
              end if;
            when q_wait5089 =>
              \$v5090\ := \$$10697_stack_ptr_take\;
              if \$v5090\(0) = '1' then
                state_var7021 <= q_wait5089;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13090_i\;
                state_var7021 <= pause_setI5087;
              end if;
            when q_wait5093 =>
              \$v5094\ := \$$10697_stack_ptr_take\;
              if \$v5094\(0) = '1' then
                state_var7021 <= q_wait5093;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5091;
              end if;
            when q_wait5097 =>
              \$v5098\ := \$$10702_brk_ptr_take\;
              if \$v5098\(0) = '1' then
                state_var7021 <= q_wait5097;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5095;
              end if;
            when q_wait5101 =>
              \$v5102\ := \$$10702_brk_ptr_take\;
              if \$v5102\(0) = '1' then
                state_var7021 <= q_wait5101;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5099;
              end if;
            when q_wait5105 =>
              \$v5106\ := \$$10702_brk_ptr_take\;
              if \$v5106\(0) = '1' then
                state_var7021 <= q_wait5105;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13098\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5103;
              end if;
            when q_wait5109 =>
              \$v5110\ := \$$10702_brk_ptr_take\;
              if \$v5110\(0) = '1' then
                state_var7021 <= q_wait5109;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5107;
              end if;
            when q_wait5114 =>
              \$v5115\ := \$$10695_limit_ptr_take\;
              if \$v5115\(0) = '1' then
                state_var7021 <= q_wait5114;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5112;
              end if;
            when q_wait5118 =>
              \$v5119\ := \$$10702_brk_ptr_take\;
              if \$v5119\(0) = '1' then
                state_var7021 <= q_wait5118;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5116;
              end if;
            when q_wait5129 =>
              \$v5130\ := \$$10697_stack_ptr_take\;
              if \$v5130\(0) = '1' then
                state_var7021 <= q_wait5129;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13084\;
                state_var7021 <= pause_setI5127;
              end if;
            when q_wait5136 =>
              \$v5137\ := \$$10696_ram_ptr_take\;
              if \$v5137\(0) = '1' then
                state_var7021 <= q_wait5136;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13079\));
                state_var7021 <= pause_getI5134;
              end if;
            when q_wait5140 =>
              \$v5141\ := \$$10697_stack_ptr_take\;
              if \$v5141\(0) = '1' then
                state_var7021 <= q_wait5140;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5138;
              end if;
            when q_wait5144 =>
              \$v5145\ := \$$10697_stack_ptr_take\;
              if \$v5145\(0) = '1' then
                state_var7021 <= q_wait5144;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13076\;
                state_var7021 <= pause_setI5142;
              end if;
            when q_wait5151 =>
              \$v5152\ := \$$10696_ram_ptr_take\;
              if \$v5152\(0) = '1' then
                state_var7021 <= q_wait5151;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13071\));
                state_var7021 <= pause_getI5149;
              end if;
            when q_wait5155 =>
              \$v5156\ := \$$10697_stack_ptr_take\;
              if \$v5156\(0) = '1' then
                state_var7021 <= q_wait5155;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5153;
              end if;
            when q_wait5160 =>
              \$v5161\ := \$$10696_ram_ptr_take\;
              if \$v5161\(0) = '1' then
                state_var7021 <= q_wait5160;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5157\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13181\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13174\ & "0000" & \$13179\ & "0001" & \$v5157\;
                state_var7021 <= pause_setI5158;
              end if;
            when q_wait5164 =>
              \$v5165\ := \$$10697_stack_ptr_take\;
              if \$v5165\(0) = '1' then
                state_var7021 <= q_wait5164;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5162;
              end if;
            when q_wait5168 =>
              \$v5169\ := \$$10697_stack_ptr_take\;
              if \$v5169\(0) = '1' then
                state_var7021 <= q_wait5168;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13178_i\;
                state_var7021 <= pause_setI5166;
              end if;
            when q_wait5172 =>
              \$v5173\ := \$$10697_stack_ptr_take\;
              if \$v5173\(0) = '1' then
                state_var7021 <= q_wait5172;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5170;
              end if;
            when q_wait5176 =>
              \$v5177\ := \$$10702_brk_ptr_take\;
              if \$v5177\(0) = '1' then
                state_var7021 <= q_wait5176;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5174;
              end if;
            when q_wait5180 =>
              \$v5181\ := \$$10702_brk_ptr_take\;
              if \$v5181\(0) = '1' then
                state_var7021 <= q_wait5180;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5178;
              end if;
            when q_wait5184 =>
              \$v5185\ := \$$10702_brk_ptr_take\;
              if \$v5185\(0) = '1' then
                state_var7021 <= q_wait5184;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13186\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5182;
              end if;
            when q_wait5188 =>
              \$v5189\ := \$$10702_brk_ptr_take\;
              if \$v5189\(0) = '1' then
                state_var7021 <= q_wait5188;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5186;
              end if;
            when q_wait5193 =>
              \$v5194\ := \$$10695_limit_ptr_take\;
              if \$v5194\(0) = '1' then
                state_var7021 <= q_wait5193;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5191;
              end if;
            when q_wait5197 =>
              \$v5198\ := \$$10702_brk_ptr_take\;
              if \$v5198\(0) = '1' then
                state_var7021 <= q_wait5197;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5195;
              end if;
            when q_wait5202 =>
              \$v5203\ := \$$10696_ram_ptr_take\;
              if \$v5203\(0) = '1' then
                state_var7021 <= q_wait5202;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5199\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13229\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13222\ & "0000" & \$13227\ & "0001" & \$v5199\;
                state_var7021 <= pause_setI5200;
              end if;
            when q_wait5206 =>
              \$v5207\ := \$$10697_stack_ptr_take\;
              if \$v5207\(0) = '1' then
                state_var7021 <= q_wait5206;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5204;
              end if;
            when q_wait5210 =>
              \$v5211\ := \$$10697_stack_ptr_take\;
              if \$v5211\(0) = '1' then
                state_var7021 <= q_wait5210;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13226_i\;
                state_var7021 <= pause_setI5208;
              end if;
            when q_wait5214 =>
              \$v5215\ := \$$10697_stack_ptr_take\;
              if \$v5215\(0) = '1' then
                state_var7021 <= q_wait5214;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5212;
              end if;
            when q_wait5218 =>
              \$v5219\ := \$$10702_brk_ptr_take\;
              if \$v5219\(0) = '1' then
                state_var7021 <= q_wait5218;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5216;
              end if;
            when q_wait5222 =>
              \$v5223\ := \$$10702_brk_ptr_take\;
              if \$v5223\(0) = '1' then
                state_var7021 <= q_wait5222;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5220;
              end if;
            when q_wait5226 =>
              \$v5227\ := \$$10702_brk_ptr_take\;
              if \$v5227\(0) = '1' then
                state_var7021 <= q_wait5226;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13234\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5224;
              end if;
            when q_wait5230 =>
              \$v5231\ := \$$10702_brk_ptr_take\;
              if \$v5231\(0) = '1' then
                state_var7021 <= q_wait5230;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5228;
              end if;
            when q_wait5235 =>
              \$v5236\ := \$$10695_limit_ptr_take\;
              if \$v5236\(0) = '1' then
                state_var7021 <= q_wait5235;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5233;
              end if;
            when q_wait5239 =>
              \$v5240\ := \$$10702_brk_ptr_take\;
              if \$v5240\(0) = '1' then
                state_var7021 <= q_wait5239;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5237;
              end if;
            when q_wait5246 =>
              \$v5247\ := \$$10697_stack_ptr_take\;
              if \$v5247\(0) = '1' then
                state_var7021 <= q_wait5246;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13220\;
                state_var7021 <= pause_setI5244;
              end if;
            when q_wait5253 =>
              \$v5254\ := \$$10696_ram_ptr_take\;
              if \$v5254\(0) = '1' then
                state_var7021 <= q_wait5253;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13215\));
                state_var7021 <= pause_getI5251;
              end if;
            when q_wait5257 =>
              \$v5258\ := \$$10697_stack_ptr_take\;
              if \$v5258\(0) = '1' then
                state_var7021 <= q_wait5257;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5255;
              end if;
            when q_wait5265 =>
              \$v5266\ := \$$10696_ram_ptr_take\;
              if \$v5266\(0) = '1' then
                state_var7021 <= q_wait5265;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13291_i\));
                state_var7021 <= pause_getI5263;
              end if;
            when q_wait5273 =>
              \$v5274\ := \$$10696_ram_ptr_take\;
              if \$v5274\(0) = '1' then
                state_var7021 <= q_wait5273;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13313_i\));
                state_var7021 <= pause_getI5271;
              end if;
            when q_wait5280 =>
              \$v5281\ := \$$10696_ram_ptr_take\;
              if \$v5281\(0) = '1' then
                state_var7021 <= q_wait5280;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13347_i\));
                state_var7021 <= pause_getI5278;
              end if;
            when q_wait5287 =>
              \$v5288\ := \$$10697_stack_ptr_take\;
              if \$v5288\(0) = '1' then
                state_var7021 <= q_wait5287;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5285;
              end if;
            when q_wait5292 =>
              \$v5293\ := \$$10696_ram_ptr_take\;
              if \$v5293\(0) = '1' then
                state_var7021 <= q_wait5292;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13368_i\));
                state_var7021 <= pause_getI5290;
              end if;
            when q_wait5301 =>
              \$v5302\ := \$$10696_ram_ptr_take\;
              if \$v5302\(0) = '1' then
                state_var7021 <= q_wait5301;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13382_i\));
                state_var7021 <= pause_getI5299;
              end if;
            when q_wait5307 =>
              \$v5308\ := \$$10700_pc_ptr_take\;
              if \$v5308\(0) = '1' then
                state_var7021 <= q_wait5307;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5305;
              end if;
            when q_wait5312 =>
              \$v5313\ := \$$10702_brk_ptr_take\;
              if \$v5313\(0) = '1' then
                state_var7021 <= q_wait5312;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5310;
              end if;
            when q_wait5316 =>
              \$v5317\ := \$$10695_limit_ptr_take\;
              if \$v5317\(0) = '1' then
                state_var7021 <= q_wait5316;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5314;
              end if;
            when q_wait5320 =>
              \$v5321\ := \$$10700_pc_ptr_take\;
              if \$v5321\(0) = '1' then
                state_var7021 <= q_wait5320;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$13415\;
                state_var7021 <= pause_setI5318;
              end if;
            when q_wait5328 =>
              \$v5329\ := \$$10696_ram_ptr_take\;
              if \$v5329\(0) = '1' then
                state_var7021 <= q_wait5328;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13442_i\));
                state_var7021 <= pause_getI5326;
              end if;
            when q_wait5334 =>
              \$v5335\ := \$$10700_pc_ptr_take\;
              if \$v5335\(0) = '1' then
                state_var7021 <= q_wait5334;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5332;
              end if;
            when q_wait5340 =>
              \$v5341\ := \$$10696_ram_ptr_take\;
              if \$v5341\(0) = '1' then
                state_var7021 <= q_wait5340;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13459_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13405\ & \$13460\(36 to 71) & \$13461\(72 to 107);
                state_var7021 <= pause_setI5338;
              end if;
            when q_wait5345 =>
              \$v5346\ := \$$10696_ram_ptr_take\;
              if \$v5346\(0) = '1' then
                state_var7021 <= q_wait5345;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13482_i\));
                state_var7021 <= pause_getI5343;
              end if;
            when q_wait5352 =>
              \$v5353\ := \$$10696_ram_ptr_take\;
              if \$v5353\(0) = '1' then
                state_var7021 <= q_wait5352;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13495_i\));
                state_var7021 <= pause_getI5350;
              end if;
            when q_wait5361 =>
              \$v5362\ := \$$10696_ram_ptr_take\;
              if \$v5362\(0) = '1' then
                state_var7021 <= q_wait5361;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13529_i\));
                state_var7021 <= pause_getI5359;
              end if;
            when q_wait5368 =>
              \$v5369\ := \$$10697_stack_ptr_take\;
              if \$v5369\(0) = '1' then
                state_var7021 <= q_wait5368;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5366;
              end if;
            when q_wait5373 =>
              \$v5374\ := \$$10696_ram_ptr_take\;
              if \$v5374\(0) = '1' then
                state_var7021 <= q_wait5373;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13545_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13405\ & \$13546\(36 to 71) & \$13547\(72 to 107);
                state_var7021 <= pause_setI5371;
              end if;
            when q_wait5378 =>
              \$v5379\ := \$$10696_ram_ptr_take\;
              if \$v5379\(0) = '1' then
                state_var7021 <= q_wait5378;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13568_i\));
                state_var7021 <= pause_getI5376;
              end if;
            when q_wait5385 =>
              \$v5386\ := \$$10696_ram_ptr_take\;
              if \$v5386\(0) = '1' then
                state_var7021 <= q_wait5385;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13581_i\));
                state_var7021 <= pause_getI5383;
              end if;
            when q_wait5395 =>
              \$v5396\ := \$$10697_stack_ptr_take\;
              if \$v5396\(0) = '1' then
                state_var7021 <= q_wait5395;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13404\;
                state_var7021 <= pause_setI5393;
              end if;
            when q_wait5402 =>
              \$v5403\ := \$$10696_ram_ptr_take\;
              if \$v5403\(0) = '1' then
                state_var7021 <= q_wait5402;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13399\));
                state_var7021 <= pause_getI5400;
              end if;
            when q_wait5406 =>
              \$v5407\ := \$$10697_stack_ptr_take\;
              if \$v5407\(0) = '1' then
                state_var7021 <= q_wait5406;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5404;
              end if;
            when q_wait5410 =>
              \$v5411\ := \$$10700_pc_ptr_take\;
              if \$v5411\(0) = '1' then
                state_var7021 <= q_wait5410;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$13613\;
                state_var7021 <= pause_setI5408;
              end if;
            when q_wait5418 =>
              \$v5419\ := \$$10696_ram_ptr_take\;
              if \$v5419\(0) = '1' then
                state_var7021 <= q_wait5418;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13640_i\));
                state_var7021 <= pause_getI5416;
              end if;
            when q_wait5424 =>
              \$v5425\ := \$$10700_pc_ptr_take\;
              if \$v5425\(0) = '1' then
                state_var7021 <= q_wait5424;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5422;
              end if;
            when q_wait5429 =>
              \$v5430\ := \$$10696_ram_ptr_take\;
              if \$v5430\(0) = '1' then
                state_var7021 <= q_wait5429;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5426\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13603\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$13596_v\ & "0000" & \$13601\ & "0001" & \$v5426\;
                state_var7021 <= pause_setI5427;
              end if;
            when q_wait5433 =>
              \$v5434\ := \$$10697_stack_ptr_take\;
              if \$v5434\(0) = '1' then
                state_var7021 <= q_wait5433;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5431;
              end if;
            when q_wait5437 =>
              \$v5438\ := \$$10697_stack_ptr_take\;
              if \$v5438\(0) = '1' then
                state_var7021 <= q_wait5437;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13600_i\;
                state_var7021 <= pause_setI5435;
              end if;
            when q_wait5441 =>
              \$v5442\ := \$$10697_stack_ptr_take\;
              if \$v5442\(0) = '1' then
                state_var7021 <= q_wait5441;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5439;
              end if;
            when q_wait5445 =>
              \$v5446\ := \$$10702_brk_ptr_take\;
              if \$v5446\(0) = '1' then
                state_var7021 <= q_wait5445;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5443;
              end if;
            when q_wait5449 =>
              \$v5450\ := \$$10702_brk_ptr_take\;
              if \$v5450\(0) = '1' then
                state_var7021 <= q_wait5449;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5447;
              end if;
            when q_wait5453 =>
              \$v5454\ := \$$10702_brk_ptr_take\;
              if \$v5454\(0) = '1' then
                state_var7021 <= q_wait5453;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13645\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5451;
              end if;
            when q_wait5457 =>
              \$v5458\ := \$$10702_brk_ptr_take\;
              if \$v5458\(0) = '1' then
                state_var7021 <= q_wait5457;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5455;
              end if;
            when q_wait5462 =>
              \$v5463\ := \$$10695_limit_ptr_take\;
              if \$v5463\(0) = '1' then
                state_var7021 <= q_wait5462;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5460;
              end if;
            when q_wait5466 =>
              \$v5467\ := \$$10702_brk_ptr_take\;
              if \$v5467\(0) = '1' then
                state_var7021 <= q_wait5466;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5464;
              end if;
            when q_wait5472 =>
              \$v5473\ := \$$10696_ram_ptr_take\;
              if \$v5473\(0) = '1' then
                state_var7021 <= q_wait5472;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13684_i\));
                state_var7021 <= pause_getI5470;
              end if;
            when q_wait5479 =>
              \$v5480\ := \$$10696_ram_ptr_take\;
              if \$v5480\(0) = '1' then
                state_var7021 <= q_wait5479;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13718_i\));
                state_var7021 <= pause_getI5477;
              end if;
            when q_wait5486 =>
              \$v5487\ := \$$10697_stack_ptr_take\;
              if \$v5487\(0) = '1' then
                state_var7021 <= q_wait5486;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5484;
              end if;
            when q_wait5491 =>
              \$v5492\ := \$$10696_ram_ptr_take\;
              if \$v5492\(0) = '1' then
                state_var7021 <= q_wait5491;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13739_i\));
                state_var7021 <= pause_getI5489;
              end if;
            when q_wait5499 =>
              \$v5500\ := \$$10700_pc_ptr_take\;
              if \$v5500\(0) = '1' then
                state_var7021 <= q_wait5499;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$13756\;
                state_var7021 <= pause_setI5497;
              end if;
            when q_wait5507 =>
              \$v5508\ := \$$10696_ram_ptr_take\;
              if \$v5508\(0) = '1' then
                state_var7021 <= q_wait5507;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13783_i\));
                state_var7021 <= pause_getI5505;
              end if;
            when q_wait5513 =>
              \$v5514\ := \$$10700_pc_ptr_take\;
              if \$v5514\(0) = '1' then
                state_var7021 <= q_wait5513;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5511;
              end if;
            when q_wait5518 =>
              \$v5519\ := \$$10696_ram_ptr_take\;
              if \$v5519\(0) = '1' then
                state_var7021 <= q_wait5518;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5515\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$13746\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$10793\(36 to 71) & "0000" & \$13744\ & "0001" & \$v5515\;
                state_var7021 <= pause_setI5516;
              end if;
            when q_wait5522 =>
              \$v5523\ := \$$10697_stack_ptr_take\;
              if \$v5523\(0) = '1' then
                state_var7021 <= q_wait5522;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5520;
              end if;
            when q_wait5526 =>
              \$v5527\ := \$$10697_stack_ptr_take\;
              if \$v5527\(0) = '1' then
                state_var7021 <= q_wait5526;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13743_i\;
                state_var7021 <= pause_setI5524;
              end if;
            when q_wait5530 =>
              \$v5531\ := \$$10697_stack_ptr_take\;
              if \$v5531\(0) = '1' then
                state_var7021 <= q_wait5530;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5528;
              end if;
            when q_wait5534 =>
              \$v5535\ := \$$10702_brk_ptr_take\;
              if \$v5535\(0) = '1' then
                state_var7021 <= q_wait5534;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5532;
              end if;
            when q_wait5538 =>
              \$v5539\ := \$$10702_brk_ptr_take\;
              if \$v5539\(0) = '1' then
                state_var7021 <= q_wait5538;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5536;
              end if;
            when q_wait5542 =>
              \$v5543\ := \$$10702_brk_ptr_take\;
              if \$v5543\(0) = '1' then
                state_var7021 <= q_wait5542;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13788\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5540;
              end if;
            when q_wait5546 =>
              \$v5547\ := \$$10702_brk_ptr_take\;
              if \$v5547\(0) = '1' then
                state_var7021 <= q_wait5546;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5544;
              end if;
            when q_wait5551 =>
              \$v5552\ := \$$10695_limit_ptr_take\;
              if \$v5552\(0) = '1' then
                state_var7021 <= q_wait5551;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5549;
              end if;
            when q_wait5555 =>
              \$v5556\ := \$$10702_brk_ptr_take\;
              if \$v5556\(0) = '1' then
                state_var7021 <= q_wait5555;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5553;
              end if;
            when q_wait5559 =>
              \$v5560\ := \$$10700_pc_ptr_take\;
              if \$v5560\(0) = '1' then
                state_var7021 <= q_wait5559;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$13837\;
                state_var7021 <= pause_setI5557;
              end if;
            when q_wait5567 =>
              \$v5568\ := \$$10696_ram_ptr_take\;
              if \$v5568\(0) = '1' then
                state_var7021 <= q_wait5567;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13864_i\));
                state_var7021 <= pause_getI5565;
              end if;
            when q_wait5573 =>
              \$v5574\ := \$$10700_pc_ptr_take\;
              if \$v5574\(0) = '1' then
                state_var7021 <= q_wait5573;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5571;
              end if;
            when q_wait5577 =>
              \$v5578\ := \$$10700_pc_ptr_take\;
              if \$v5578\(0) = '1' then
                state_var7021 <= q_wait5577;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$13816\;
                state_var7021 <= pause_setI5575;
              end if;
            when q_wait5596 =>
              \$v5597\ := \$$10697_stack_ptr_take\;
              if \$v5597\(0) = '1' then
                state_var7021 <= q_wait5596;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$13812\;
                state_var7021 <= pause_setI5594;
              end if;
            when q_wait5603 =>
              \$v5604\ := \$$10696_ram_ptr_take\;
              if \$v5604\(0) = '1' then
                state_var7021 <= q_wait5603;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13807\));
                state_var7021 <= pause_getI5601;
              end if;
            when q_wait5607 =>
              \$v5608\ := \$$10697_stack_ptr_take\;
              if \$v5608\(0) = '1' then
                state_var7021 <= q_wait5607;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI5605;
              end if;
            when q_wait5615 =>
              \$v5616\ := \$$10696_ram_ptr_take\;
              if \$v5616\(0) = '1' then
                state_var7021 <= q_wait5615;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13913_i\));
                state_var7021 <= pause_getI5613;
              end if;
            when q_wait5621 =>
              \$v5622\ := \$$10700_pc_ptr_take\;
              if \$v5622\(0) = '1' then
                state_var7021 <= q_wait5621;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr\ <= 0;
                state_var7021 <= pause_getI5619;
              end if;
            when q_wait5625 =>
              \$v5626\ := \$$10697_stack_ptr_take\;
              if \$v5626\(0) = '1' then
                state_var7021 <= q_wait5625;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$10767_j\;
                state_var7021 <= pause_setI5623;
              end if;
            when q_wait5631 =>
              \$v5632\ := \$$10696_ram_ptr_take\;
              if \$v5632\(0) = '1' then
                state_var7021 <= q_wait5631;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5627\ := X"0000000" & X"0";
                \$v5628\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10767_j\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5627\ & "0001" & \$v5628\ & "0000" & \$10763_i\;
                state_var7021 <= pause_setI5629;
              end if;
            when q_wait5638 =>
              \$v5639\ := \$$10696_ram_ptr_take\;
              if \$v5639\(0) = '1' then
                state_var7021 <= q_wait5638;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5633\ := X"0000000" & X"5";
                \$v5634\ := X"0000000" & X"0";
                \$v5635\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$10763_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5633\ & "0001" & \$v5634\ & "0001" & \$v5635\;
                state_var7021 <= pause_setI5636;
              end if;
            when q_wait5642 =>
              \$v5643\ := \$$10702_brk_ptr_take\;
              if \$v5643\(0) = '1' then
                state_var7021 <= q_wait5642;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5640;
              end if;
            when q_wait5646 =>
              \$v5647\ := \$$10702_brk_ptr_take\;
              if \$v5647\(0) = '1' then
                state_var7021 <= q_wait5646;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5644;
              end if;
            when q_wait5650 =>
              \$v5651\ := \$$10702_brk_ptr_take\;
              if \$v5651\(0) = '1' then
                state_var7021 <= q_wait5650;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13923\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5648;
              end if;
            when q_wait5654 =>
              \$v5655\ := \$$10702_brk_ptr_take\;
              if \$v5655\(0) = '1' then
                state_var7021 <= q_wait5654;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5652;
              end if;
            when q_wait5659 =>
              \$v5660\ := \$$10695_limit_ptr_take\;
              if \$v5660\(0) = '1' then
                state_var7021 <= q_wait5659;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5657;
              end if;
            when q_wait5663 =>
              \$v5664\ := \$$10702_brk_ptr_take\;
              if \$v5664\(0) = '1' then
                state_var7021 <= q_wait5663;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5661;
              end if;
            when q_wait5667 =>
              \$v5668\ := \$$10702_brk_ptr_take\;
              if \$v5668\(0) = '1' then
                state_var7021 <= q_wait5667;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5665;
              end if;
            when q_wait5671 =>
              \$v5672\ := \$$10702_brk_ptr_take\;
              if \$v5672\(0) = '1' then
                state_var7021 <= q_wait5671;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5669;
              end if;
            when q_wait5675 =>
              \$v5676\ := \$$10702_brk_ptr_take\;
              if \$v5676\(0) = '1' then
                state_var7021 <= q_wait5675;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$13942\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5673;
              end if;
            when q_wait5679 =>
              \$v5680\ := \$$10702_brk_ptr_take\;
              if \$v5680\(0) = '1' then
                state_var7021 <= q_wait5679;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5677;
              end if;
            when q_wait5684 =>
              \$v5685\ := \$$10695_limit_ptr_take\;
              if \$v5685\(0) = '1' then
                state_var7021 <= q_wait5684;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5682;
              end if;
            when q_wait5688 =>
              \$v5689\ := \$$10702_brk_ptr_take\;
              if \$v5689\(0) = '1' then
                state_var7021 <= q_wait5688;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5686;
              end if;
            when q_wait5692 =>
              \$v5693\ := \$$10699_symtbl_ptr_take\;
              if \$v5693\(0) = '1' then
                state_var7021 <= q_wait5692;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$13972\;
                state_var7021 <= pause_setI5690;
              end if;
            when q_wait5700 =>
              \$v5701\ := \$$10696_ram_ptr_take\;
              if \$v5701\(0) = '1' then
                state_var7021 <= q_wait5700;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$13999_i\));
                state_var7021 <= pause_getI5698;
              end if;
            when q_wait5706 =>
              \$v5707\ := \$$10699_symtbl_ptr_take\;
              if \$v5707\(0) = '1' then
                state_var7021 <= q_wait5706;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5704;
              end if;
            when q_wait5712 =>
              \$v5713\ := \$$10696_ram_ptr_take\;
              if \$v5713\(0) = '1' then
                state_var7021 <= q_wait5712;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5709\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14012_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v5709\ & \$14017\(36 to 71) & \$14022\(72 to 107);
                state_var7021 <= pause_setI5710;
              end if;
            when q_wait5717 =>
              \$v5718\ := \$$10696_ram_ptr_take\;
              if \$v5718\(0) = '1' then
                state_var7021 <= q_wait5717;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14045_i\));
                state_var7021 <= pause_getI5715;
              end if;
            when q_wait5724 =>
              \$v5725\ := \$$10696_ram_ptr_take\;
              if \$v5725\(0) = '1' then
                state_var7021 <= q_wait5724;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14058_i\));
                state_var7021 <= pause_getI5722;
              end if;
            when q_wait5733 =>
              \$v5734\ := \$$10696_ram_ptr_take\;
              if \$v5734\(0) = '1' then
                state_var7021 <= q_wait5733;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14072_i\));
                state_var7021 <= pause_getI5731;
              end if;
            when q_wait5739 =>
              \$v5740\ := \$$10699_symtbl_ptr_take\;
              if \$v5740\(0) = '1' then
                state_var7021 <= q_wait5739;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5737;
              end if;
            when q_wait5743 =>
              \$v5744\ := \$$10699_symtbl_ptr_take\;
              if \$v5744\(0) = '1' then
                state_var7021 <= q_wait5743;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$14085\;
                state_var7021 <= pause_setI5741;
              end if;
            when q_wait5751 =>
              \$v5752\ := \$$10696_ram_ptr_take\;
              if \$v5752\(0) = '1' then
                state_var7021 <= q_wait5751;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14112_i\));
                state_var7021 <= pause_getI5749;
              end if;
            when q_wait5757 =>
              \$v5758\ := \$$10699_symtbl_ptr_take\;
              if \$v5758\(0) = '1' then
                state_var7021 <= q_wait5757;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5755;
              end if;
            when q_wait5763 =>
              \$v5764\ := \$$10696_ram_ptr_take\;
              if \$v5764\(0) = '1' then
                state_var7021 <= q_wait5763;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5760\ := X"0000000" & X"1";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14125_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v5760\ & \$14130\(36 to 71) & \$14135\(72 to 107);
                state_var7021 <= pause_setI5761;
              end if;
            when q_wait5768 =>
              \$v5769\ := \$$10696_ram_ptr_take\;
              if \$v5769\(0) = '1' then
                state_var7021 <= q_wait5768;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14158_i\));
                state_var7021 <= pause_getI5766;
              end if;
            when q_wait5775 =>
              \$v5776\ := \$$10696_ram_ptr_take\;
              if \$v5776\(0) = '1' then
                state_var7021 <= q_wait5775;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14171_i\));
                state_var7021 <= pause_getI5773;
              end if;
            when q_wait5784 =>
              \$v5785\ := \$$10696_ram_ptr_take\;
              if \$v5785\(0) = '1' then
                state_var7021 <= q_wait5784;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14185_i\));
                state_var7021 <= pause_getI5782;
              end if;
            when q_wait5790 =>
              \$v5791\ := \$$10699_symtbl_ptr_take\;
              if \$v5791\(0) = '1' then
                state_var7021 <= q_wait5790;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5788;
              end if;
            when q_wait5794 =>
              \$v5795\ := \$$10699_symtbl_ptr_take\;
              if \$v5795\(0) = '1' then
                state_var7021 <= q_wait5794;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$14198\;
                state_var7021 <= pause_setI5792;
              end if;
            when q_wait5802 =>
              \$v5803\ := \$$10696_ram_ptr_take\;
              if \$v5803\(0) = '1' then
                state_var7021 <= q_wait5802;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14225_i\));
                state_var7021 <= pause_getI5800;
              end if;
            when q_wait5808 =>
              \$v5809\ := \$$10699_symtbl_ptr_take\;
              if \$v5809\(0) = '1' then
                state_var7021 <= q_wait5808;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5806;
              end if;
            when q_wait5814 =>
              \$v5815\ := \$$10696_ram_ptr_take\;
              if \$v5815\(0) = '1' then
                state_var7021 <= q_wait5814;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5811\ := X"0000000" & X"2";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14238_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v5811\ & \$14243\(36 to 71) & \$14248\(72 to 107);
                state_var7021 <= pause_setI5812;
              end if;
            when q_wait5819 =>
              \$v5820\ := \$$10696_ram_ptr_take\;
              if \$v5820\(0) = '1' then
                state_var7021 <= q_wait5819;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14271_i\));
                state_var7021 <= pause_getI5817;
              end if;
            when q_wait5826 =>
              \$v5827\ := \$$10696_ram_ptr_take\;
              if \$v5827\(0) = '1' then
                state_var7021 <= q_wait5826;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14284_i\));
                state_var7021 <= pause_getI5824;
              end if;
            when q_wait5835 =>
              \$v5836\ := \$$10696_ram_ptr_take\;
              if \$v5836\(0) = '1' then
                state_var7021 <= q_wait5835;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14298_i\));
                state_var7021 <= pause_getI5833;
              end if;
            when q_wait5841 =>
              \$v5842\ := \$$10699_symtbl_ptr_take\;
              if \$v5842\(0) = '1' then
                state_var7021 <= q_wait5841;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5839;
              end if;
            when q_wait5845 =>
              \$v5846\ := \$$10699_symtbl_ptr_take\;
              if \$v5846\(0) = '1' then
                state_var7021 <= q_wait5845;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$14306\;
                state_var7021 <= pause_setI5843;
              end if;
            when q_wait5853 =>
              \$v5854\ := \$$10696_ram_ptr_take\;
              if \$v5854\(0) = '1' then
                state_var7021 <= q_wait5853;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14333_i\));
                state_var7021 <= pause_getI5851;
              end if;
            when q_wait5859 =>
              \$v5860\ := \$$10699_symtbl_ptr_take\;
              if \$v5860\(0) = '1' then
                state_var7021 <= q_wait5859;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5857;
              end if;
            when q_wait5864 =>
              \$v5865\ := \$$10696_ram_ptr_take\;
              if \$v5865\(0) = '1' then
                state_var7021 <= q_wait5864;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14346_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$10738_main_rib\ & \$14351\(36 to 71) & \$14356\(72 to 107);
                state_var7021 <= pause_setI5862;
              end if;
            when q_wait5869 =>
              \$v5870\ := \$$10696_ram_ptr_take\;
              if \$v5870\(0) = '1' then
                state_var7021 <= q_wait5869;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14377_i\));
                state_var7021 <= pause_getI5867;
              end if;
            when q_wait5876 =>
              \$v5877\ := \$$10696_ram_ptr_take\;
              if \$v5877\(0) = '1' then
                state_var7021 <= q_wait5876;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14390_i\));
                state_var7021 <= pause_getI5874;
              end if;
            when q_wait5885 =>
              \$v5886\ := \$$10696_ram_ptr_take\;
              if \$v5886\(0) = '1' then
                state_var7021 <= q_wait5885;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14404_i\));
                state_var7021 <= pause_getI5883;
              end if;
            when q_wait5891 =>
              \$v5892\ := \$$10699_symtbl_ptr_take\;
              if \$v5892\(0) = '1' then
                state_var7021 <= q_wait5891;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5889;
              end if;
            when q_wait5895 =>
              \$v5896\ := \$$10698_heap_ptr_take\;
              if \$v5896\(0) = '1' then
                state_var7021 <= q_wait5895;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5893;
              end if;
            when q_wait5901 =>
              \$v5902\ := \$$10696_ram_ptr_take\;
              if \$v5902\(0) = '1' then
                state_var7021 <= q_wait5901;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5897\ := X"0000000" & X"0";
                \$v5898\ := X"0000000" & X"1";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14407\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5897\ & "0000" & \$10734\ & "0001" & \$v5898\;
                state_var7021 <= pause_setI5899;
              end if;
            when q_wait5905 =>
              \$v5906\ := \$$10698_heap_ptr_take\;
              if \$v5906\(0) = '1' then
                state_var7021 <= q_wait5905;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5903;
              end if;
            when q_wait5909 =>
              \$v5910\ := \$$10698_heap_ptr_take\;
              if \$v5910\(0) = '1' then
                state_var7021 <= q_wait5909;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14405_i\;
                state_var7021 <= pause_setI5907;
              end if;
            when q_wait5913 =>
              \$v5914\ := \$$10702_brk_ptr_take\;
              if \$v5914\(0) = '1' then
                state_var7021 <= q_wait5913;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5911;
              end if;
            when q_wait5917 =>
              \$v5918\ := \$$10702_brk_ptr_take\;
              if \$v5918\(0) = '1' then
                state_var7021 <= q_wait5917;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5915;
              end if;
            when q_wait5921 =>
              \$v5922\ := \$$10702_brk_ptr_take\;
              if \$v5922\(0) = '1' then
                state_var7021 <= q_wait5921;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14415\ & X"0000000" & X"1");
                state_var7021 <= pause_setI5919;
              end if;
            when q_wait5925 =>
              \$v5926\ := \$$10702_brk_ptr_take\;
              if \$v5926\(0) = '1' then
                state_var7021 <= q_wait5925;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5923;
              end if;
            when q_wait5930 =>
              \$v5931\ := \$$10695_limit_ptr_take\;
              if \$v5931\(0) = '1' then
                state_var7021 <= q_wait5930;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI5928;
              end if;
            when q_wait5934 =>
              \$v5935\ := \$$10702_brk_ptr_take\;
              if \$v5935\(0) = '1' then
                state_var7021 <= q_wait5934;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI5932;
              end if;
            when q_wait5938 =>
              \$v5939\ := \$$10699_symtbl_ptr_take\;
              if \$v5939\(0) = '1' then
                state_var7021 <= q_wait5938;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI5936;
              end if;
            when q_wait5942 =>
              \$v5943\ := \$$10700_pc_ptr_take\;
              if \$v5943\(0) = '1' then
                state_var7021 <= q_wait5942;
              else
                \$$10700_pc_ptr_take\(0) := '1';
                \$$10700_pc_ptr_write\ <= 0;
                \$$10700_pc_write_request\ <= '1';
                \$$10700_pc_write\ <= \$10731\;
                state_var7021 <= pause_setI5940;
              end if;
            when q_wait5950 =>
              \$v5951\ := \$$10696_ram_ptr_take\;
              if \$v5951\(0) = '1' then
                state_var7021 <= q_wait5950;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14458_i\));
                state_var7021 <= pause_getI5948;
              end if;
            when q_wait5957 =>
              \$v5958\ := \$$10696_ram_ptr_take\;
              if \$v5958\(0) = '1' then
                state_var7021 <= q_wait5957;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14472_i\));
                state_var7021 <= pause_getI5955;
              end if;
            when q_wait5963 =>
              \$v5964\ := \$$10698_heap_ptr_take\;
              if \$v5964\(0) = '1' then
                state_var7021 <= q_wait5963;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5961;
              end if;
            when q_wait5968 =>
              \$v5969\ := \$$10696_ram_ptr_take\;
              if \$v5969\(0) = '1' then
                state_var7021 <= q_wait5968;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15090_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15076_new_rib\ & \$15091\(36 to 71) & \$15092\(72 to 107);
                state_var7021 <= pause_setI5966;
              end if;
            when q_wait5973 =>
              \$v5974\ := \$$10696_ram_ptr_take\;
              if \$v5974\(0) = '1' then
                state_var7021 <= q_wait5973;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15114_i\));
                state_var7021 <= pause_getI5971;
              end if;
            when q_wait5980 =>
              \$v5981\ := \$$10696_ram_ptr_take\;
              if \$v5981\(0) = '1' then
                state_var7021 <= q_wait5980;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15128_i\));
                state_var7021 <= pause_getI5978;
              end if;
            when q_wait5988 =>
              \$v5989\ := \$$10698_heap_ptr_take\;
              if \$v5989\(0) = '1' then
                state_var7021 <= q_wait5988;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5986;
              end if;
            when q_wait5993 =>
              \$v5994\ := \$$10696_ram_ptr_take\;
              if \$v5994\(0) = '1' then
                state_var7021 <= q_wait5993;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v5990\ := X"0000000" & X"4";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15131\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v5990\ & \$15068_opnd\ & \$15071\(0 to 35);
                state_var7021 <= pause_setI5991;
              end if;
            when q_wait5997 =>
              \$v5998\ := \$$10698_heap_ptr_take\;
              if \$v5998\(0) = '1' then
                state_var7021 <= q_wait5997;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI5995;
              end if;
            when q_wait6001 =>
              \$v6002\ := \$$10698_heap_ptr_take\;
              if \$v6002\(0) = '1' then
                state_var7021 <= q_wait6001;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$15129_i\;
                state_var7021 <= pause_setI5999;
              end if;
            when q_wait6005 =>
              \$v6006\ := \$$10702_brk_ptr_take\;
              if \$v6006\(0) = '1' then
                state_var7021 <= q_wait6005;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6003;
              end if;
            when q_wait6009 =>
              \$v6010\ := \$$10702_brk_ptr_take\;
              if \$v6010\(0) = '1' then
                state_var7021 <= q_wait6009;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6007;
              end if;
            when q_wait6013 =>
              \$v6014\ := \$$10702_brk_ptr_take\;
              if \$v6014\(0) = '1' then
                state_var7021 <= q_wait6013;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15141\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6011;
              end if;
            when q_wait6017 =>
              \$v6018\ := \$$10702_brk_ptr_take\;
              if \$v6018\(0) = '1' then
                state_var7021 <= q_wait6017;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6015;
              end if;
            when q_wait6022 =>
              \$v6023\ := \$$10695_limit_ptr_take\;
              if \$v6023\(0) = '1' then
                state_var7021 <= q_wait6022;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6020;
              end if;
            when q_wait6026 =>
              \$v6027\ := \$$10702_brk_ptr_take\;
              if \$v6027\(0) = '1' then
                state_var7021 <= q_wait6026;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6024;
              end if;
            when q_wait6031 =>
              \$v6032\ := \$$10696_ram_ptr_take\;
              if \$v6032\(0) = '1' then
                state_var7021 <= q_wait6031;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15172_i\));
                state_var7021 <= pause_getI6029;
              end if;
            when q_wait6037 =>
              \$v6038\ := \$$10697_stack_ptr_take\;
              if \$v6038\(0) = '1' then
                state_var7021 <= q_wait6037;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6035;
              end if;
            when q_wait6041 =>
              \$v6042\ := \$$10697_stack_ptr_take\;
              if \$v6042\(0) = '1' then
                state_var7021 <= q_wait6041;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$15067\;
                state_var7021 <= pause_setI6039;
              end if;
            when q_wait6048 =>
              \$v6049\ := \$$10696_ram_ptr_take\;
              if \$v6049\(0) = '1' then
                state_var7021 <= q_wait6048;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15062\));
                state_var7021 <= pause_getI6046;
              end if;
            when q_wait6052 =>
              \$v6053\ := \$$10697_stack_ptr_take\;
              if \$v6053\(0) = '1' then
                state_var7021 <= q_wait6052;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6050;
              end if;
            when q_wait6057 =>
              \$v6058\ := \$$10696_ram_ptr_take\;
              if \$v6058\(0) = '1' then
                state_var7021 <= q_wait6057;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14681_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$14667_new_rib\ & \$14682\(36 to 71) & \$14683\(72 to 107);
                state_var7021 <= pause_setI6055;
              end if;
            when q_wait6062 =>
              \$v6063\ := \$$10696_ram_ptr_take\;
              if \$v6063\(0) = '1' then
                state_var7021 <= q_wait6062;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14705_i\));
                state_var7021 <= pause_getI6060;
              end if;
            when q_wait6069 =>
              \$v6070\ := \$$10696_ram_ptr_take\;
              if \$v6070\(0) = '1' then
                state_var7021 <= q_wait6069;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14719_i\));
                state_var7021 <= pause_getI6067;
              end if;
            when q_wait6077 =>
              \$v6078\ := \$$10698_heap_ptr_take\;
              if \$v6078\(0) = '1' then
                state_var7021 <= q_wait6077;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6075;
              end if;
            when q_wait6082 =>
              \$v6083\ := \$$10696_ram_ptr_take\;
              if \$v6083\(0) = '1' then
                state_var7021 <= q_wait6082;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6079\ := X"0000000" & X"3";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14722\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v6079\ & \$14656_proc_rib\ & \$14662\(0 to 35);
                state_var7021 <= pause_setI6080;
              end if;
            when q_wait6086 =>
              \$v6087\ := \$$10698_heap_ptr_take\;
              if \$v6087\(0) = '1' then
                state_var7021 <= q_wait6086;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6084;
              end if;
            when q_wait6090 =>
              \$v6091\ := \$$10698_heap_ptr_take\;
              if \$v6091\(0) = '1' then
                state_var7021 <= q_wait6090;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14720_i\;
                state_var7021 <= pause_setI6088;
              end if;
            when q_wait6094 =>
              \$v6095\ := \$$10702_brk_ptr_take\;
              if \$v6095\(0) = '1' then
                state_var7021 <= q_wait6094;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6092;
              end if;
            when q_wait6098 =>
              \$v6099\ := \$$10702_brk_ptr_take\;
              if \$v6099\(0) = '1' then
                state_var7021 <= q_wait6098;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6096;
              end if;
            when q_wait6102 =>
              \$v6103\ := \$$10702_brk_ptr_take\;
              if \$v6103\(0) = '1' then
                state_var7021 <= q_wait6102;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14732\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6100;
              end if;
            when q_wait6106 =>
              \$v6107\ := \$$10702_brk_ptr_take\;
              if \$v6107\(0) = '1' then
                state_var7021 <= q_wait6106;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6104;
              end if;
            when q_wait6111 =>
              \$v6112\ := \$$10695_limit_ptr_take\;
              if \$v6112\(0) = '1' then
                state_var7021 <= q_wait6111;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6109;
              end if;
            when q_wait6115 =>
              \$v6116\ := \$$10702_brk_ptr_take\;
              if \$v6116\(0) = '1' then
                state_var7021 <= q_wait6115;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6113;
              end if;
            when q_wait6120 =>
              \$v6121\ := \$$10696_ram_ptr_take\;
              if \$v6121\(0) = '1' then
                state_var7021 <= q_wait6120;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14763_i\));
                state_var7021 <= pause_getI6118;
              end if;
            when q_wait6126 =>
              \$v6127\ := \$$10697_stack_ptr_take\;
              if \$v6127\(0) = '1' then
                state_var7021 <= q_wait6126;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6124;
              end if;
            when q_wait6134 =>
              \$v6135\ := \$$10697_stack_ptr_take\;
              if \$v6135\(0) = '1' then
                state_var7021 <= q_wait6134;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6132;
              end if;
            when q_wait6138 =>
              \$v6139\ := \$$10698_heap_ptr_take\;
              if \$v6139\(0) = '1' then
                state_var7021 <= q_wait6138;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6136;
              end if;
            when q_wait6144 =>
              \$v6145\ := \$$10696_ram_ptr_take\;
              if \$v6145\(0) = '1' then
                state_var7021 <= q_wait6144;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6140\ := X"0000000" & X"0";
                \$v6141\ := X"0000000" & X"1";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14770\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$14652_code_proc_rib\ & "0000" & \$v6140\ & "0001" & \$v6141\;
                state_var7021 <= pause_setI6142;
              end if;
            when q_wait6148 =>
              \$v6149\ := \$$10698_heap_ptr_take\;
              if \$v6149\(0) = '1' then
                state_var7021 <= q_wait6148;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6146;
              end if;
            when q_wait6152 =>
              \$v6153\ := \$$10698_heap_ptr_take\;
              if \$v6153\(0) = '1' then
                state_var7021 <= q_wait6152;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14768_i\;
                state_var7021 <= pause_setI6150;
              end if;
            when q_wait6156 =>
              \$v6157\ := \$$10702_brk_ptr_take\;
              if \$v6157\(0) = '1' then
                state_var7021 <= q_wait6156;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6154;
              end if;
            when q_wait6160 =>
              \$v6161\ := \$$10702_brk_ptr_take\;
              if \$v6161\(0) = '1' then
                state_var7021 <= q_wait6160;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6158;
              end if;
            when q_wait6164 =>
              \$v6165\ := \$$10702_brk_ptr_take\;
              if \$v6165\(0) = '1' then
                state_var7021 <= q_wait6164;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14777\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6162;
              end if;
            when q_wait6168 =>
              \$v6169\ := \$$10702_brk_ptr_take\;
              if \$v6169\(0) = '1' then
                state_var7021 <= q_wait6168;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6166;
              end if;
            when q_wait6173 =>
              \$v6174\ := \$$10695_limit_ptr_take\;
              if \$v6174\(0) = '1' then
                state_var7021 <= q_wait6173;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6171;
              end if;
            when q_wait6177 =>
              \$v6178\ := \$$10702_brk_ptr_take\;
              if \$v6178\(0) = '1' then
                state_var7021 <= q_wait6177;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6175;
              end if;
            when q_wait6181 =>
              \$v6182\ := \$$10698_heap_ptr_take\;
              if \$v6182\(0) = '1' then
                state_var7021 <= q_wait6181;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6179;
              end if;
            when q_wait6186 =>
              \$v6187\ := \$$10696_ram_ptr_take\;
              if \$v6187\(0) = '1' then
                state_var7021 <= q_wait6186;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6183\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14797\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$14533_opnd\ & "0001" & \$v6183\ & \$14648_ty\;
                state_var7021 <= pause_setI6184;
              end if;
            when q_wait6190 =>
              \$v6191\ := \$$10698_heap_ptr_take\;
              if \$v6191\(0) = '1' then
                state_var7021 <= q_wait6190;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6188;
              end if;
            when q_wait6194 =>
              \$v6195\ := \$$10698_heap_ptr_take\;
              if \$v6195\(0) = '1' then
                state_var7021 <= q_wait6194;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14795_i\;
                state_var7021 <= pause_setI6192;
              end if;
            when q_wait6198 =>
              \$v6199\ := \$$10702_brk_ptr_take\;
              if \$v6199\(0) = '1' then
                state_var7021 <= q_wait6198;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6196;
              end if;
            when q_wait6202 =>
              \$v6203\ := \$$10702_brk_ptr_take\;
              if \$v6203\(0) = '1' then
                state_var7021 <= q_wait6202;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6200;
              end if;
            when q_wait6206 =>
              \$v6207\ := \$$10702_brk_ptr_take\;
              if \$v6207\(0) = '1' then
                state_var7021 <= q_wait6206;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14803\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6204;
              end if;
            when q_wait6210 =>
              \$v6211\ := \$$10702_brk_ptr_take\;
              if \$v6211\(0) = '1' then
                state_var7021 <= q_wait6210;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6208;
              end if;
            when q_wait6215 =>
              \$v6216\ := \$$10695_limit_ptr_take\;
              if \$v6216\(0) = '1' then
                state_var7021 <= q_wait6215;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6213;
              end if;
            when q_wait6219 =>
              \$v6220\ := \$$10702_brk_ptr_take\;
              if \$v6220\(0) = '1' then
                state_var7021 <= q_wait6219;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6217;
              end if;
            when q_wait6223 =>
              \$v6224\ := \$$10697_stack_ptr_take\;
              if \$v6224\(0) = '1' then
                state_var7021 <= q_wait6223;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$14647\;
                state_var7021 <= pause_setI6221;
              end if;
            when q_wait6230 =>
              \$v6231\ := \$$10696_ram_ptr_take\;
              if \$v6231\(0) = '1' then
                state_var7021 <= q_wait6230;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14642\));
                state_var7021 <= pause_getI6228;
              end if;
            when q_wait6234 =>
              \$v6235\ := \$$10697_stack_ptr_take\;
              if \$v6235\(0) = '1' then
                state_var7021 <= q_wait6234;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6232;
              end if;
            when q_wait6239 =>
              \$v6240\ := \$$10696_ram_ptr_take\;
              if \$v6240\(0) = '1' then
                state_var7021 <= q_wait6239;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14556_i\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$14542_new_rib\ & \$14557\(36 to 71) & \$14558\(72 to 107);
                state_var7021 <= pause_setI6237;
              end if;
            when q_wait6244 =>
              \$v6245\ := \$$10696_ram_ptr_take\;
              if \$v6245\(0) = '1' then
                state_var7021 <= q_wait6244;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14580_i\));
                state_var7021 <= pause_getI6242;
              end if;
            when q_wait6251 =>
              \$v6252\ := \$$10696_ram_ptr_take\;
              if \$v6252\(0) = '1' then
                state_var7021 <= q_wait6251;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14594_i\));
                state_var7021 <= pause_getI6249;
              end if;
            when q_wait6259 =>
              \$v6260\ := \$$10698_heap_ptr_take\;
              if \$v6260\(0) = '1' then
                state_var7021 <= q_wait6259;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6257;
              end if;
            when q_wait6264 =>
              \$v6265\ := \$$10696_ram_ptr_take\;
              if \$v6265\(0) = '1' then
                state_var7021 <= q_wait6264;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6261\ := eclat_if(eclat_lt(X"0000000" & X"0" & \$14511_loop311_arg\(0 to 31)) & eclat_sub(\$14511_loop311_arg\(0 to 31) & X"0000000" & X"1") & X"0000000" & X"0");
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$14597\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v6261\ & \$14533_opnd\ & \$14537\(0 to 35);
                state_var7021 <= pause_setI6262;
              end if;
            when q_wait6268 =>
              \$v6269\ := \$$10698_heap_ptr_take\;
              if \$v6269\(0) = '1' then
                state_var7021 <= q_wait6268;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6266;
              end if;
            when q_wait6272 =>
              \$v6273\ := \$$10698_heap_ptr_take\;
              if \$v6273\(0) = '1' then
                state_var7021 <= q_wait6272;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$14595_i\;
                state_var7021 <= pause_setI6270;
              end if;
            when q_wait6276 =>
              \$v6277\ := \$$10702_brk_ptr_take\;
              if \$v6277\(0) = '1' then
                state_var7021 <= q_wait6276;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6274;
              end if;
            when q_wait6280 =>
              \$v6281\ := \$$10702_brk_ptr_take\;
              if \$v6281\(0) = '1' then
                state_var7021 <= q_wait6280;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6278;
              end if;
            when q_wait6284 =>
              \$v6285\ := \$$10702_brk_ptr_take\;
              if \$v6285\(0) = '1' then
                state_var7021 <= q_wait6284;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$14609\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6282;
              end if;
            when q_wait6288 =>
              \$v6289\ := \$$10702_brk_ptr_take\;
              if \$v6289\(0) = '1' then
                state_var7021 <= q_wait6288;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6286;
              end if;
            when q_wait6293 =>
              \$v6294\ := \$$10695_limit_ptr_take\;
              if \$v6294\(0) = '1' then
                state_var7021 <= q_wait6293;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6291;
              end if;
            when q_wait6297 =>
              \$v6298\ := \$$10702_brk_ptr_take\;
              if \$v6298\(0) = '1' then
                state_var7021 <= q_wait6297;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6295;
              end if;
            when q_wait6302 =>
              \$v6303\ := \$$10696_ram_ptr_take\;
              if \$v6303\(0) = '1' then
                state_var7021 <= q_wait6302;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14640_i\));
                state_var7021 <= pause_getI6300;
              end if;
            when q_wait6308 =>
              \$v6309\ := \$$10697_stack_ptr_take\;
              if \$v6309\(0) = '1' then
                state_var7021 <= q_wait6308;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6306;
              end if;
            when q_wait6314 =>
              \$v6315\ := \$$10696_ram_ptr_take\;
              if \$v6315\(0) = '1' then
                state_var7021 <= q_wait6314;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14991_i\));
                state_var7021 <= pause_getI6312;
              end if;
            when q_wait6321 =>
              \$v6322\ := \$$10696_ram_ptr_take\;
              if \$v6322\(0) = '1' then
                state_var7021 <= q_wait6321;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15025_i\));
                state_var7021 <= pause_getI6319;
              end if;
            when q_wait6328 =>
              \$v6329\ := \$$10699_symtbl_ptr_take\;
              if \$v6329\(0) = '1' then
                state_var7021 <= q_wait6328;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6326;
              end if;
            when q_wait6335 =>
              \$v6336\ := \$$10701_pos_ptr_take\;
              if \$v6336\(0) = '1' then
                state_var7021 <= q_wait6335;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$14948\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6333;
              end if;
            when q_wait6339 =>
              \$v6340\ := \$$10701_pos_ptr_take\;
              if \$v6340\(0) = '1' then
                state_var7021 <= q_wait6339;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6337;
              end if;
            when q_wait6343 =>
              \$v6344\ := \$$10701_pos_ptr_take\;
              if \$v6344\(0) = '1' then
                state_var7021 <= q_wait6343;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6341;
              end if;
            when q_wait6348 =>
              \$v6349\ := \$$10696_ram_ptr_take\;
              if \$v6349\(0) = '1' then
                state_var7021 <= q_wait6348;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14858_i\));
                state_var7021 <= pause_getI6346;
              end if;
            when q_wait6355 =>
              \$v6356\ := \$$10696_ram_ptr_take\;
              if \$v6356\(0) = '1' then
                state_var7021 <= q_wait6355;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$14892_i\));
                state_var7021 <= pause_getI6353;
              end if;
            when q_wait6362 =>
              \$v6363\ := \$$10699_symtbl_ptr_take\;
              if \$v6363\(0) = '1' then
                state_var7021 <= q_wait6362;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6360;
              end if;
            when q_wait6367 =>
              \$v6368\ := \$$10701_pos_ptr_take\;
              if \$v6368\(0) = '1' then
                state_var7021 <= q_wait6367;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$14912\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6365;
              end if;
            when q_wait6371 =>
              \$v6372\ := \$$10701_pos_ptr_take\;
              if \$v6372\(0) = '1' then
                state_var7021 <= q_wait6371;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6369;
              end if;
            when q_wait6375 =>
              \$v6376\ := \$$10701_pos_ptr_take\;
              if \$v6376\(0) = '1' then
                state_var7021 <= q_wait6375;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6373;
              end if;
            when q_wait6383 =>
              \$v6384\ := \$$10696_ram_ptr_take\;
              if \$v6384\(0) = '1' then
                state_var7021 <= q_wait6383;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6379\ := \$14511_loop311_arg\(0 to 31);
                \$v6380\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15037\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v6379\ & "0000" & \$15035\ & "0001" & \$v6380\;
                state_var7021 <= pause_setI6381;
              end if;
            when q_wait6387 =>
              \$v6388\ := \$$10697_stack_ptr_take\;
              if \$v6388\(0) = '1' then
                state_var7021 <= q_wait6387;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6385;
              end if;
            when q_wait6391 =>
              \$v6392\ := \$$10697_stack_ptr_take\;
              if \$v6392\(0) = '1' then
                state_var7021 <= q_wait6391;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= \$15034_i\;
                state_var7021 <= pause_setI6389;
              end if;
            when q_wait6395 =>
              \$v6396\ := \$$10697_stack_ptr_take\;
              if \$v6396\(0) = '1' then
                state_var7021 <= q_wait6395;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr\ <= 0;
                state_var7021 <= pause_getI6393;
              end if;
            when q_wait6399 =>
              \$v6400\ := \$$10702_brk_ptr_take\;
              if \$v6400\(0) = '1' then
                state_var7021 <= q_wait6399;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6397;
              end if;
            when q_wait6403 =>
              \$v6404\ := \$$10702_brk_ptr_take\;
              if \$v6404\(0) = '1' then
                state_var7021 <= q_wait6403;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6401;
              end if;
            when q_wait6407 =>
              \$v6408\ := \$$10702_brk_ptr_take\;
              if \$v6408\(0) = '1' then
                state_var7021 <= q_wait6407;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15043\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6405;
              end if;
            when q_wait6411 =>
              \$v6412\ := \$$10702_brk_ptr_take\;
              if \$v6412\(0) = '1' then
                state_var7021 <= q_wait6411;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6409;
              end if;
            when q_wait6416 =>
              \$v6417\ := \$$10695_limit_ptr_take\;
              if \$v6417\(0) = '1' then
                state_var7021 <= q_wait6416;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6414;
              end if;
            when q_wait6420 =>
              \$v6421\ := \$$10702_brk_ptr_take\;
              if \$v6421\(0) = '1' then
                state_var7021 <= q_wait6420;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6418;
              end if;
            when q_wait6427 =>
              \$v6428\ := \$$10701_pos_ptr_take\;
              if \$v6428\(0) = '1' then
                state_var7021 <= q_wait6427;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$14499\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6425;
              end if;
            when q_wait6431 =>
              \$v6432\ := \$$10701_pos_ptr_take\;
              if \$v6432\(0) = '1' then
                state_var7021 <= q_wait6431;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6429;
              end if;
            when q_wait6435 =>
              \$v6436\ := \$$10701_pos_ptr_take\;
              if \$v6436\(0) = '1' then
                state_var7021 <= q_wait6435;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6433;
              end if;
            when q_wait6439 =>
              \$v6440\ := \$$10699_symtbl_ptr_take\;
              if \$v6440\(0) = '1' then
                state_var7021 <= q_wait6439;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6437;
              end if;
            when q_wait6444 =>
              \$v6445\ := \$$10696_ram_ptr_take\;
              if \$v6445\(0) = '1' then
                state_var7021 <= q_wait6444;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6441\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15648\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15642_end_rib\ & "0000" & \$15621\ & "0001" & \$v6441\;
                state_var7021 <= pause_setI6442;
              end if;
            when q_wait6448 =>
              \$v6449\ := \$$10699_symtbl_ptr_take\;
              if \$v6449\(0) = '1' then
                state_var7021 <= q_wait6448;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6446;
              end if;
            when q_wait6452 =>
              \$v6453\ := \$$10699_symtbl_ptr_take\;
              if \$v6453\(0) = '1' then
                state_var7021 <= q_wait6452;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15646_i\;
                state_var7021 <= pause_setI6450;
              end if;
            when q_wait6456 =>
              \$v6457\ := \$$10702_brk_ptr_take\;
              if \$v6457\(0) = '1' then
                state_var7021 <= q_wait6456;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6454;
              end if;
            when q_wait6460 =>
              \$v6461\ := \$$10702_brk_ptr_take\;
              if \$v6461\(0) = '1' then
                state_var7021 <= q_wait6460;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6458;
              end if;
            when q_wait6464 =>
              \$v6465\ := \$$10702_brk_ptr_take\;
              if \$v6465\(0) = '1' then
                state_var7021 <= q_wait6464;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15655\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6462;
              end if;
            when q_wait6468 =>
              \$v6469\ := \$$10702_brk_ptr_take\;
              if \$v6469\(0) = '1' then
                state_var7021 <= q_wait6468;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6466;
              end if;
            when q_wait6473 =>
              \$v6474\ := \$$10695_limit_ptr_take\;
              if \$v6474\(0) = '1' then
                state_var7021 <= q_wait6473;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6471;
              end if;
            when q_wait6477 =>
              \$v6478\ := \$$10702_brk_ptr_take\;
              if \$v6478\(0) = '1' then
                state_var7021 <= q_wait6477;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6475;
              end if;
            when q_wait6481 =>
              \$v6482\ := \$$10699_symtbl_ptr_take\;
              if \$v6482\(0) = '1' then
                state_var7021 <= q_wait6481;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6479;
              end if;
            when q_wait6487 =>
              \$v6488\ := \$$10696_ram_ptr_take\;
              if \$v6488\(0) = '1' then
                state_var7021 <= q_wait6487;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6483\ := X"0000000" & X"2";
                \$v6484\ := X"0000000" & X"2";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15640\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v6483\ & \$15634_str_rib\ & "0001" & \$v6484\;
                state_var7021 <= pause_setI6485;
              end if;
            when q_wait6491 =>
              \$v6492\ := \$$10699_symtbl_ptr_take\;
              if \$v6492\(0) = '1' then
                state_var7021 <= q_wait6491;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6489;
              end if;
            when q_wait6495 =>
              \$v6496\ := \$$10699_symtbl_ptr_take\;
              if \$v6496\(0) = '1' then
                state_var7021 <= q_wait6495;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15638_i\;
                state_var7021 <= pause_setI6493;
              end if;
            when q_wait6499 =>
              \$v6500\ := \$$10702_brk_ptr_take\;
              if \$v6500\(0) = '1' then
                state_var7021 <= q_wait6499;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6497;
              end if;
            when q_wait6503 =>
              \$v6504\ := \$$10702_brk_ptr_take\;
              if \$v6504\(0) = '1' then
                state_var7021 <= q_wait6503;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6501;
              end if;
            when q_wait6507 =>
              \$v6508\ := \$$10702_brk_ptr_take\;
              if \$v6508\(0) = '1' then
                state_var7021 <= q_wait6507;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15678\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6505;
              end if;
            when q_wait6511 =>
              \$v6512\ := \$$10702_brk_ptr_take\;
              if \$v6512\(0) = '1' then
                state_var7021 <= q_wait6511;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6509;
              end if;
            when q_wait6516 =>
              \$v6517\ := \$$10695_limit_ptr_take\;
              if \$v6517\(0) = '1' then
                state_var7021 <= q_wait6516;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6514;
              end if;
            when q_wait6520 =>
              \$v6521\ := \$$10702_brk_ptr_take\;
              if \$v6521\(0) = '1' then
                state_var7021 <= q_wait6520;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6518;
              end if;
            when q_wait6524 =>
              \$v6525\ := \$$10699_symtbl_ptr_take\;
              if \$v6525\(0) = '1' then
                state_var7021 <= q_wait6524;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6522;
              end if;
            when q_wait6530 =>
              \$v6531\ := \$$10696_ram_ptr_take\;
              if \$v6531\(0) = '1' then
                state_var7021 <= q_wait6530;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6526\ := X"0000000" & X"0";
                \$v6527\ := X"0000000" & X"3";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15632\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v6526\ & "0001" & \$15622\ & "0001" & \$v6527\;
                state_var7021 <= pause_setI6528;
              end if;
            when q_wait6534 =>
              \$v6535\ := \$$10699_symtbl_ptr_take\;
              if \$v6535\(0) = '1' then
                state_var7021 <= q_wait6534;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6532;
              end if;
            when q_wait6538 =>
              \$v6539\ := \$$10699_symtbl_ptr_take\;
              if \$v6539\(0) = '1' then
                state_var7021 <= q_wait6538;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15630_i\;
                state_var7021 <= pause_setI6536;
              end if;
            when q_wait6542 =>
              \$v6543\ := \$$10702_brk_ptr_take\;
              if \$v6543\(0) = '1' then
                state_var7021 <= q_wait6542;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6540;
              end if;
            when q_wait6546 =>
              \$v6547\ := \$$10702_brk_ptr_take\;
              if \$v6547\(0) = '1' then
                state_var7021 <= q_wait6546;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6544;
              end if;
            when q_wait6550 =>
              \$v6551\ := \$$10702_brk_ptr_take\;
              if \$v6551\(0) = '1' then
                state_var7021 <= q_wait6550;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15702\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6548;
              end if;
            when q_wait6554 =>
              \$v6555\ := \$$10702_brk_ptr_take\;
              if \$v6555\(0) = '1' then
                state_var7021 <= q_wait6554;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6552;
              end if;
            when q_wait6559 =>
              \$v6560\ := \$$10695_limit_ptr_take\;
              if \$v6560\(0) = '1' then
                state_var7021 <= q_wait6559;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6557;
              end if;
            when q_wait6563 =>
              \$v6564\ := \$$10702_brk_ptr_take\;
              if \$v6564\(0) = '1' then
                state_var7021 <= q_wait6563;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6561;
              end if;
            when q_wait6568 =>
              \$v6569\ := \$$10696_ram_ptr_take\;
              if \$v6569\(0) = '1' then
                state_var7021 <= q_wait6568;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15754_i\));
                state_var7021 <= pause_getI6566;
              end if;
            when q_wait6587 =>
              \$v6588\ := \$$10696_ram_ptr_take\;
              if \$v6588\(0) = '1' then
                state_var7021 <= q_wait6587;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15780_i\));
                state_var7021 <= pause_getI6585;
              end if;
            when q_wait6598 =>
              \$v6599\ := \$$10699_symtbl_ptr_take\;
              if \$v6599\(0) = '1' then
                state_var7021 <= q_wait6598;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6596;
              end if;
            when q_wait6603 =>
              \$v6604\ := \$$10699_symtbl_ptr_take\;
              if \$v6604\(0) = '1' then
                state_var7021 <= q_wait6603;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6601;
              end if;
            when q_wait6608 =>
              \$v6609\ := \$$10696_ram_ptr_take\;
              if \$v6609\(0) = '1' then
                state_var7021 <= q_wait6608;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6605\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15481\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15475_end_rib\ & "0000" & \$15454\ & "0001" & \$v6605\;
                state_var7021 <= pause_setI6606;
              end if;
            when q_wait6612 =>
              \$v6613\ := \$$10699_symtbl_ptr_take\;
              if \$v6613\(0) = '1' then
                state_var7021 <= q_wait6612;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6610;
              end if;
            when q_wait6616 =>
              \$v6617\ := \$$10699_symtbl_ptr_take\;
              if \$v6617\(0) = '1' then
                state_var7021 <= q_wait6616;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15479_i\;
                state_var7021 <= pause_setI6614;
              end if;
            when q_wait6620 =>
              \$v6621\ := \$$10702_brk_ptr_take\;
              if \$v6621\(0) = '1' then
                state_var7021 <= q_wait6620;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6618;
              end if;
            when q_wait6624 =>
              \$v6625\ := \$$10702_brk_ptr_take\;
              if \$v6625\(0) = '1' then
                state_var7021 <= q_wait6624;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6622;
              end if;
            when q_wait6628 =>
              \$v6629\ := \$$10702_brk_ptr_take\;
              if \$v6629\(0) = '1' then
                state_var7021 <= q_wait6628;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15488\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6626;
              end if;
            when q_wait6632 =>
              \$v6633\ := \$$10702_brk_ptr_take\;
              if \$v6633\(0) = '1' then
                state_var7021 <= q_wait6632;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6630;
              end if;
            when q_wait6637 =>
              \$v6638\ := \$$10695_limit_ptr_take\;
              if \$v6638\(0) = '1' then
                state_var7021 <= q_wait6637;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6635;
              end if;
            when q_wait6641 =>
              \$v6642\ := \$$10702_brk_ptr_take\;
              if \$v6642\(0) = '1' then
                state_var7021 <= q_wait6641;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6639;
              end if;
            when q_wait6645 =>
              \$v6646\ := \$$10699_symtbl_ptr_take\;
              if \$v6646\(0) = '1' then
                state_var7021 <= q_wait6645;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6643;
              end if;
            when q_wait6651 =>
              \$v6652\ := \$$10696_ram_ptr_take\;
              if \$v6652\(0) = '1' then
                state_var7021 <= q_wait6651;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6647\ := X"0000000" & X"2";
                \$v6648\ := X"0000000" & X"2";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15473\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v6647\ & \$15467_str_rib\ & "0001" & \$v6648\;
                state_var7021 <= pause_setI6649;
              end if;
            when q_wait6655 =>
              \$v6656\ := \$$10699_symtbl_ptr_take\;
              if \$v6656\(0) = '1' then
                state_var7021 <= q_wait6655;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6653;
              end if;
            when q_wait6659 =>
              \$v6660\ := \$$10699_symtbl_ptr_take\;
              if \$v6660\(0) = '1' then
                state_var7021 <= q_wait6659;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15471_i\;
                state_var7021 <= pause_setI6657;
              end if;
            when q_wait6663 =>
              \$v6664\ := \$$10702_brk_ptr_take\;
              if \$v6664\(0) = '1' then
                state_var7021 <= q_wait6663;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6661;
              end if;
            when q_wait6667 =>
              \$v6668\ := \$$10702_brk_ptr_take\;
              if \$v6668\(0) = '1' then
                state_var7021 <= q_wait6667;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6665;
              end if;
            when q_wait6671 =>
              \$v6672\ := \$$10702_brk_ptr_take\;
              if \$v6672\(0) = '1' then
                state_var7021 <= q_wait6671;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15511\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6669;
              end if;
            when q_wait6675 =>
              \$v6676\ := \$$10702_brk_ptr_take\;
              if \$v6676\(0) = '1' then
                state_var7021 <= q_wait6675;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6673;
              end if;
            when q_wait6680 =>
              \$v6681\ := \$$10695_limit_ptr_take\;
              if \$v6681\(0) = '1' then
                state_var7021 <= q_wait6680;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6678;
              end if;
            when q_wait6684 =>
              \$v6685\ := \$$10702_brk_ptr_take\;
              if \$v6685\(0) = '1' then
                state_var7021 <= q_wait6684;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6682;
              end if;
            when q_wait6688 =>
              \$v6689\ := \$$10699_symtbl_ptr_take\;
              if \$v6689\(0) = '1' then
                state_var7021 <= q_wait6688;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6686;
              end if;
            when q_wait6693 =>
              \$v6694\ := \$$10696_ram_ptr_take\;
              if \$v6694\(0) = '1' then
                state_var7021 <= q_wait6693;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6690\ := X"0000000" & X"3";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15465\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15240_loop23133355_arg\(0 to 35) & "0001" & \$15455\ & "0001" & \$v6690\;
                state_var7021 <= pause_setI6691;
              end if;
            when q_wait6697 =>
              \$v6698\ := \$$10699_symtbl_ptr_take\;
              if \$v6698\(0) = '1' then
                state_var7021 <= q_wait6697;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6695;
              end if;
            when q_wait6701 =>
              \$v6702\ := \$$10699_symtbl_ptr_take\;
              if \$v6702\(0) = '1' then
                state_var7021 <= q_wait6701;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15463_i\;
                state_var7021 <= pause_setI6699;
              end if;
            when q_wait6705 =>
              \$v6706\ := \$$10702_brk_ptr_take\;
              if \$v6706\(0) = '1' then
                state_var7021 <= q_wait6705;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6703;
              end if;
            when q_wait6709 =>
              \$v6710\ := \$$10702_brk_ptr_take\;
              if \$v6710\(0) = '1' then
                state_var7021 <= q_wait6709;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6707;
              end if;
            when q_wait6713 =>
              \$v6714\ := \$$10702_brk_ptr_take\;
              if \$v6714\(0) = '1' then
                state_var7021 <= q_wait6713;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15534\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6711;
              end if;
            when q_wait6717 =>
              \$v6718\ := \$$10702_brk_ptr_take\;
              if \$v6718\(0) = '1' then
                state_var7021 <= q_wait6717;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6715;
              end if;
            when q_wait6722 =>
              \$v6723\ := \$$10695_limit_ptr_take\;
              if \$v6723\(0) = '1' then
                state_var7021 <= q_wait6722;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6720;
              end if;
            when q_wait6726 =>
              \$v6727\ := \$$10702_brk_ptr_take\;
              if \$v6727\(0) = '1' then
                state_var7021 <= q_wait6726;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6724;
              end if;
            when q_wait6731 =>
              \$v6732\ := \$$10696_ram_ptr_take\;
              if \$v6732\(0) = '1' then
                state_var7021 <= q_wait6731;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15585_i\));
                state_var7021 <= pause_getI6729;
              end if;
            when q_wait6750 =>
              \$v6751\ := \$$10696_ram_ptr_take\;
              if \$v6751\(0) = '1' then
                state_var7021 <= q_wait6750;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15611_i\));
                state_var7021 <= pause_getI6748;
              end if;
            when q_wait6760 =>
              \$v6761\ := \$$10699_symtbl_ptr_take\;
              if \$v6761\(0) = '1' then
                state_var7021 <= q_wait6760;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6758;
              end if;
            when q_wait6764 =>
              \$v6765\ := \$$10699_symtbl_ptr_take\;
              if \$v6765\(0) = '1' then
                state_var7021 <= q_wait6764;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6762;
              end if;
            when q_wait6769 =>
              \$v6770\ := \$$10696_ram_ptr_take\;
              if \$v6770\(0) = '1' then
                state_var7021 <= q_wait6769;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6766\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15317\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15311_end_rib\ & "0000" & \$15293\ & "0001" & \$v6766\;
                state_var7021 <= pause_setI6767;
              end if;
            when q_wait6773 =>
              \$v6774\ := \$$10699_symtbl_ptr_take\;
              if \$v6774\(0) = '1' then
                state_var7021 <= q_wait6773;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6771;
              end if;
            when q_wait6777 =>
              \$v6778\ := \$$10699_symtbl_ptr_take\;
              if \$v6778\(0) = '1' then
                state_var7021 <= q_wait6777;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15315_i\;
                state_var7021 <= pause_setI6775;
              end if;
            when q_wait6781 =>
              \$v6782\ := \$$10702_brk_ptr_take\;
              if \$v6782\(0) = '1' then
                state_var7021 <= q_wait6781;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6779;
              end if;
            when q_wait6785 =>
              \$v6786\ := \$$10702_brk_ptr_take\;
              if \$v6786\(0) = '1' then
                state_var7021 <= q_wait6785;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6783;
              end if;
            when q_wait6789 =>
              \$v6790\ := \$$10702_brk_ptr_take\;
              if \$v6790\(0) = '1' then
                state_var7021 <= q_wait6789;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15324\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6787;
              end if;
            when q_wait6793 =>
              \$v6794\ := \$$10702_brk_ptr_take\;
              if \$v6794\(0) = '1' then
                state_var7021 <= q_wait6793;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6791;
              end if;
            when q_wait6798 =>
              \$v6799\ := \$$10695_limit_ptr_take\;
              if \$v6799\(0) = '1' then
                state_var7021 <= q_wait6798;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6796;
              end if;
            when q_wait6802 =>
              \$v6803\ := \$$10702_brk_ptr_take\;
              if \$v6803\(0) = '1' then
                state_var7021 <= q_wait6802;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6800;
              end if;
            when q_wait6806 =>
              \$v6807\ := \$$10699_symtbl_ptr_take\;
              if \$v6807\(0) = '1' then
                state_var7021 <= q_wait6806;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6804;
              end if;
            when q_wait6812 =>
              \$v6813\ := \$$10696_ram_ptr_take\;
              if \$v6813\(0) = '1' then
                state_var7021 <= q_wait6812;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6808\ := X"0000000" & X"2";
                \$v6809\ := X"0000000" & X"2";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15309\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0000" & \$v6808\ & \$15303_str_rib\ & "0001" & \$v6809\;
                state_var7021 <= pause_setI6810;
              end if;
            when q_wait6816 =>
              \$v6817\ := \$$10699_symtbl_ptr_take\;
              if \$v6817\(0) = '1' then
                state_var7021 <= q_wait6816;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6814;
              end if;
            when q_wait6820 =>
              \$v6821\ := \$$10699_symtbl_ptr_take\;
              if \$v6821\(0) = '1' then
                state_var7021 <= q_wait6820;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15307_i\;
                state_var7021 <= pause_setI6818;
              end if;
            when q_wait6824 =>
              \$v6825\ := \$$10702_brk_ptr_take\;
              if \$v6825\(0) = '1' then
                state_var7021 <= q_wait6824;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6822;
              end if;
            when q_wait6828 =>
              \$v6829\ := \$$10702_brk_ptr_take\;
              if \$v6829\(0) = '1' then
                state_var7021 <= q_wait6828;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6826;
              end if;
            when q_wait6832 =>
              \$v6833\ := \$$10702_brk_ptr_take\;
              if \$v6833\(0) = '1' then
                state_var7021 <= q_wait6832;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15347\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6830;
              end if;
            when q_wait6836 =>
              \$v6837\ := \$$10702_brk_ptr_take\;
              if \$v6837\(0) = '1' then
                state_var7021 <= q_wait6836;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6834;
              end if;
            when q_wait6841 =>
              \$v6842\ := \$$10695_limit_ptr_take\;
              if \$v6842\(0) = '1' then
                state_var7021 <= q_wait6841;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6839;
              end if;
            when q_wait6845 =>
              \$v6846\ := \$$10702_brk_ptr_take\;
              if \$v6846\(0) = '1' then
                state_var7021 <= q_wait6845;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6843;
              end if;
            when q_wait6849 =>
              \$v6850\ := \$$10699_symtbl_ptr_take\;
              if \$v6850\(0) = '1' then
                state_var7021 <= q_wait6849;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6847;
              end if;
            when q_wait6854 =>
              \$v6855\ := \$$10696_ram_ptr_take\;
              if \$v6855\(0) = '1' then
                state_var7021 <= q_wait6854;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6851\ := X"0000000" & X"3";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15301\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= \$15240_loop23133355_arg\(0 to 35) & "0001" & \$15294\ & "0001" & \$v6851\;
                state_var7021 <= pause_setI6852;
              end if;
            when q_wait6858 =>
              \$v6859\ := \$$10699_symtbl_ptr_take\;
              if \$v6859\(0) = '1' then
                state_var7021 <= q_wait6858;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6856;
              end if;
            when q_wait6862 =>
              \$v6863\ := \$$10699_symtbl_ptr_take\;
              if \$v6863\(0) = '1' then
                state_var7021 <= q_wait6862;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= \$15299_i\;
                state_var7021 <= pause_setI6860;
              end if;
            when q_wait6866 =>
              \$v6867\ := \$$10702_brk_ptr_take\;
              if \$v6867\(0) = '1' then
                state_var7021 <= q_wait6866;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6864;
              end if;
            when q_wait6870 =>
              \$v6871\ := \$$10702_brk_ptr_take\;
              if \$v6871\(0) = '1' then
                state_var7021 <= q_wait6870;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6868;
              end if;
            when q_wait6874 =>
              \$v6875\ := \$$10702_brk_ptr_take\;
              if \$v6875\(0) = '1' then
                state_var7021 <= q_wait6874;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15370\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6872;
              end if;
            when q_wait6878 =>
              \$v6879\ := \$$10702_brk_ptr_take\;
              if \$v6879\(0) = '1' then
                state_var7021 <= q_wait6878;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6876;
              end if;
            when q_wait6883 =>
              \$v6884\ := \$$10695_limit_ptr_take\;
              if \$v6884\(0) = '1' then
                state_var7021 <= q_wait6883;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6881;
              end if;
            when q_wait6887 =>
              \$v6888\ := \$$10702_brk_ptr_take\;
              if \$v6888\(0) = '1' then
                state_var7021 <= q_wait6887;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6885;
              end if;
            when q_wait6892 =>
              \$v6893\ := \$$10696_ram_ptr_take\;
              if \$v6893\(0) = '1' then
                state_var7021 <= q_wait6892;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15421_i\));
                state_var7021 <= pause_getI6890;
              end if;
            when q_wait6911 =>
              \$v6912\ := \$$10696_ram_ptr_take\;
              if \$v6912\(0) = '1' then
                state_var7021 <= q_wait6911;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$$10696_ram_ptr\ <= to_integer(unsigned(\$15447_i\));
                state_var7021 <= pause_getI6909;
              end if;
            when q_wait6921 =>
              \$v6922\ := \$$10699_symtbl_ptr_take\;
              if \$v6922\(0) = '1' then
                state_var7021 <= q_wait6921;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr\ <= 0;
                state_var7021 <= pause_getI6919;
              end if;
            when q_wait6925 =>
              \$v6926\ := \$$10698_heap_ptr_take\;
              if \$v6926\(0) = '1' then
                state_var7021 <= q_wait6925;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6923;
              end if;
            when q_wait6931 =>
              \$v6932\ := \$$10696_ram_ptr_take\;
              if \$v6932\(0) = '1' then
                state_var7021 <= q_wait6931;
              else
                \$$10696_ram_ptr_take\(0) := '1';
                \$v6927\ := eclat_vector_get(X"000000" & X"29" & X"000000" & X"3b" & X"000000" & X"27" & X"000000" & X"75" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"44" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"41" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3a" & X"000000" & X"3f" & X"000000" & X"3e" & X"000000" & X"76" & X"000000" & X"52" & X"000000" & X"3d" & X"000000" & X"21" & X"000000" & X"28" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"6d" & X"000000" & X"21" & X"000000" & X"27" & X"000000" & X"3a" & X"000000" & X"6c" & X"000000" & X"6b" & X"000000" & X"76" & X"000000" & X"36" & X"000000" & X"79" & \$15255\,32);
                \$v6928\ := X"0000000" & X"0";
                \$$10696_ram_ptr_write\ <= to_integer(unsigned(\$15265\));
                \$$10696_ram_write_request\ <= '1';
                \$$10696_ram_write\ <= "0001" & \$v6927\ & \$15240_loop23133355_arg\(0 to 35) & "0001" & \$v6928\;
                state_var7021 <= pause_setI6929;
              end if;
            when q_wait6935 =>
              \$v6936\ := \$$10698_heap_ptr_take\;
              if \$v6936\(0) = '1' then
                state_var7021 <= q_wait6935;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr\ <= 0;
                state_var7021 <= pause_getI6933;
              end if;
            when q_wait6939 =>
              \$v6940\ := \$$10698_heap_ptr_take\;
              if \$v6940\(0) = '1' then
                state_var7021 <= q_wait6939;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= \$15263_i\;
                state_var7021 <= pause_setI6937;
              end if;
            when q_wait6943 =>
              \$v6944\ := \$$10702_brk_ptr_take\;
              if \$v6944\(0) = '1' then
                state_var7021 <= q_wait6943;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6941;
              end if;
            when q_wait6947 =>
              \$v6948\ := \$$10702_brk_ptr_take\;
              if \$v6948\(0) = '1' then
                state_var7021 <= q_wait6947;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6945;
              end if;
            when q_wait6951 =>
              \$v6952\ := \$$10702_brk_ptr_take\;
              if \$v6952\(0) = '1' then
                state_var7021 <= q_wait6951;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= eclat_add(\$15274\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6949;
              end if;
            when q_wait6955 =>
              \$v6956\ := \$$10702_brk_ptr_take\;
              if \$v6956\(0) = '1' then
                state_var7021 <= q_wait6955;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6953;
              end if;
            when q_wait6960 =>
              \$v6961\ := \$$10695_limit_ptr_take\;
              if \$v6961\(0) = '1' then
                state_var7021 <= q_wait6960;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr\ <= 0;
                state_var7021 <= pause_getI6958;
              end if;
            when q_wait6964 =>
              \$v6965\ := \$$10702_brk_ptr_take\;
              if \$v6965\(0) = '1' then
                state_var7021 <= q_wait6964;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr\ <= 0;
                state_var7021 <= pause_getI6962;
              end if;
            when q_wait6970 =>
              \$v6971\ := \$$10701_pos_ptr_take\;
              if \$v6971\(0) = '1' then
                state_var7021 <= q_wait6970;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$15256\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6968;
              end if;
            when q_wait6974 =>
              \$v6975\ := \$$10701_pos_ptr_take\;
              if \$v6975\(0) = '1' then
                state_var7021 <= q_wait6974;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6972;
              end if;
            when q_wait6978 =>
              \$v6979\ := \$$10701_pos_ptr_take\;
              if \$v6979\(0) = '1' then
                state_var7021 <= q_wait6978;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6976;
              end if;
            when q_wait6985 =>
              \$v6986\ := \$$10701_pos_ptr_take\;
              if \$v6986\(0) = '1' then
                state_var7021 <= q_wait6985;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= eclat_add(\$15797\ & X"0000000" & X"1");
                state_var7021 <= pause_setI6983;
              end if;
            when q_wait6989 =>
              \$v6990\ := \$$10701_pos_ptr_take\;
              if \$v6990\(0) = '1' then
                state_var7021 <= q_wait6989;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6987;
              end if;
            when q_wait6993 =>
              \$v6994\ := \$$10701_pos_ptr_take\;
              if \$v6994\(0) = '1' then
                state_var7021 <= q_wait6993;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr\ <= 0;
                state_var7021 <= pause_getI6991;
              end if;
            when q_wait6997 =>
              \$v6998\ := \$$10695_limit_ptr_take\;
              if \$v6998\(0) = '1' then
                state_var7021 <= q_wait6997;
              else
                \$$10695_limit_ptr_take\(0) := '1';
                \$$10695_limit_ptr_write\ <= 0;
                \$$10695_limit_write_request\ <= '1';
                \$$10695_limit_write\ <= eclat_div(X"0000" & X"2710" & X"0000000" & X"2");
                state_var7021 <= pause_setI6995;
              end if;
            when q_wait7001 =>
              \$v7002\ := \$$10702_brk_ptr_take\;
              if \$v7002\(0) = '1' then
                state_var7021 <= q_wait7001;
              else
                \$$10702_brk_ptr_take\(0) := '1';
                \$$10702_brk_ptr_write\ <= 0;
                \$$10702_brk_write_request\ <= '1';
                \$$10702_brk_write\ <= X"0000000" & X"4";
                state_var7021 <= pause_setI6999;
              end if;
            when q_wait7005 =>
              \$v7006\ := \$$10701_pos_ptr_take\;
              if \$v7006\(0) = '1' then
                state_var7021 <= q_wait7005;
              else
                \$$10701_pos_ptr_take\(0) := '1';
                \$$10701_pos_ptr_write\ <= 0;
                \$$10701_pos_write_request\ <= '1';
                \$$10701_pos_write\ <= X"0000000" & X"0";
                state_var7021 <= pause_setI7003;
              end if;
            when q_wait7009 =>
              \$v7010\ := \$$10699_symtbl_ptr_take\;
              if \$v7010\(0) = '1' then
                state_var7021 <= q_wait7009;
              else
                \$$10699_symtbl_ptr_take\(0) := '1';
                \$$10699_symtbl_ptr_write\ <= 0;
                \$$10699_symtbl_write_request\ <= '1';
                \$$10699_symtbl_write\ <= eclat_sub(X"0000000" & X"0" & X"0000000" & X"1");
                state_var7021 <= pause_setI7007;
              end if;
            when q_wait7013 =>
              \$v7014\ := \$$10698_heap_ptr_take\;
              if \$v7014\(0) = '1' then
                state_var7021 <= q_wait7013;
              else
                \$$10698_heap_ptr_take\(0) := '1';
                \$$10698_heap_ptr_write\ <= 0;
                \$$10698_heap_write_request\ <= '1';
                \$$10698_heap_write\ <= eclat_sub(X"0000000" & X"0" & X"0000000" & X"1");
                state_var7021 <= pause_setI7011;
              end if;
            when q_wait7017 =>
              \$v7018\ := \$$10697_stack_ptr_take\;
              if \$v7018\(0) = '1' then
                state_var7021 <= q_wait7017;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= eclat_sub(X"0000000" & X"0" & X"0000000" & X"1");
                state_var7021 <= pause_setI7015;
              end if;
            when compute3367 =>
              rdy3366 := eclat_false;
              eclat_print_string(of_string("RVM"));
              
              eclat_print_newline(eclat_unit);
              
              \$v7018\ := \$$10697_stack_ptr_take\;
              if \$v7018\(0) = '1' then
                state_var7021 <= q_wait7017;
              else
                \$$10697_stack_ptr_take\(0) := '1';
                \$$10697_stack_ptr_write\ <= 0;
                \$$10697_stack_write_request\ <= '1';
                \$$10697_stack_write\ <= eclat_sub(X"0000000" & X"0" & X"0000000" & X"1");
                state_var7021 <= pause_setI7015;
              end if;
            end case;
            \$v7020\ := eclat_not(rdy3366);
            if \$v7020\(0) = '1' then
              result3365 := eclat_unit;
            end if;
            result3362 := result3365 & rdy3366;
            rdy3363 := eclat_true;
            state <= compute3364;
          end case;
          
          result <= result3362;
          rdy <= rdy3363;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
